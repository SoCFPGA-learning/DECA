-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"0b0b0b0b",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"00000016",
     7 => x"00000000",
     8 => x"0b0b80c0",
     9 => x"dc080b0b",
    10 => x"80c0e008",
    11 => x"0b0b80c0",
    12 => x"e4080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b80",
    15 => x"c0e40c0b",
    16 => x"0b80c0e0",
    17 => x"0c0b0b80",
    18 => x"c0dc0c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b0bb784",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"80c0dc70",
    57 => x"80cb9827",
    58 => x"8b388071",
    59 => x"70840553",
    60 => x"0c81e304",
    61 => x"8c5189b4",
    62 => x"0402fc05",
    63 => x"0df88051",
    64 => x"8f0b80c0",
    65 => x"ec0c9f0b",
    66 => x"80c0f00c",
    67 => x"a0717081",
    68 => x"05533480",
    69 => x"c0f008ff",
    70 => x"0580c0f0",
    71 => x"0c80c0f0",
    72 => x"088025e8",
    73 => x"3880c0ec",
    74 => x"08ff0580",
    75 => x"c0ec0c80",
    76 => x"c0ec0880",
    77 => x"25d03880",
    78 => x"0b80c0f0",
    79 => x"0c800b80",
    80 => x"c0ec0c02",
    81 => x"84050d04",
    82 => x"02f0050d",
    83 => x"f88053f8",
    84 => x"a05483bf",
    85 => x"52737081",
    86 => x"05553351",
    87 => x"70737081",
    88 => x"055534ff",
    89 => x"12527180",
    90 => x"25eb38fb",
    91 => x"c0539f52",
    92 => x"a0737081",
    93 => x"055534ff",
    94 => x"12527180",
    95 => x"25f23802",
    96 => x"90050d04",
    97 => x"02f4050d",
    98 => x"74538e0b",
    99 => x"80c0ec08",
   100 => x"25913882",
   101 => x"c82d80c0",
   102 => x"ec08ff05",
   103 => x"80c0ec0c",
   104 => x"838a0480",
   105 => x"c0ec0880",
   106 => x"c0f00853",
   107 => x"51728a2e",
   108 => x"098106be",
   109 => x"38715171",
   110 => x"9f24a438",
   111 => x"80c0ec08",
   112 => x"a02911f8",
   113 => x"80115151",
   114 => x"a0713480",
   115 => x"c0f00881",
   116 => x"0580c0f0",
   117 => x"0c80c0f0",
   118 => x"08519f71",
   119 => x"25de3880",
   120 => x"0b80c0f0",
   121 => x"0c80c0ec",
   122 => x"08810580",
   123 => x"c0ec0c84",
   124 => x"880470a0",
   125 => x"2912f880",
   126 => x"11515172",
   127 => x"713480c0",
   128 => x"f0088105",
   129 => x"80c0f00c",
   130 => x"80c0f008",
   131 => x"a02e0981",
   132 => x"06913880",
   133 => x"0b80c0f0",
   134 => x"0c80c0ec",
   135 => x"08810580",
   136 => x"c0ec0c02",
   137 => x"8c050d04",
   138 => x"02e8050d",
   139 => x"77795656",
   140 => x"880bfc16",
   141 => x"77712c8f",
   142 => x"06545254",
   143 => x"80537272",
   144 => x"25953871",
   145 => x"53fbe014",
   146 => x"51877134",
   147 => x"8114ff14",
   148 => x"545472f1",
   149 => x"387153f9",
   150 => x"1576712c",
   151 => x"87065351",
   152 => x"71802e8b",
   153 => x"38fbe014",
   154 => x"51717134",
   155 => x"81145472",
   156 => x"8e249538",
   157 => x"8f733153",
   158 => x"fbe01451",
   159 => x"a0713481",
   160 => x"14ff1454",
   161 => x"5472f138",
   162 => x"0298050d",
   163 => x"0402ec05",
   164 => x"0d800b80",
   165 => x"c0f40cf6",
   166 => x"8c08f690",
   167 => x"0871882c",
   168 => x"565481ff",
   169 => x"06527372",
   170 => x"25893871",
   171 => x"54820b80",
   172 => x"c0f40c72",
   173 => x"882c7381",
   174 => x"ff065455",
   175 => x"7473258d",
   176 => x"387280c0",
   177 => x"f4088407",
   178 => x"80c0f40c",
   179 => x"5573842b",
   180 => x"86a07125",
   181 => x"83713170",
   182 => x"0b0b0bbc",
   183 => x"bc0c8171",
   184 => x"2bff05f6",
   185 => x"880cfdfc",
   186 => x"13ff122c",
   187 => x"788829ff",
   188 => x"94057081",
   189 => x"2c80c0f4",
   190 => x"08525852",
   191 => x"55515254",
   192 => x"76802e85",
   193 => x"38708107",
   194 => x"5170f694",
   195 => x"0c710981",
   196 => x"05f6800c",
   197 => x"72098105",
   198 => x"f6840c02",
   199 => x"94050d04",
   200 => x"02f4050d",
   201 => x"74537270",
   202 => x"81055480",
   203 => x"f52d5271",
   204 => x"802e8938",
   205 => x"71518384",
   206 => x"2d86a604",
   207 => x"810b80c0",
   208 => x"dc0c028c",
   209 => x"050d0402",
   210 => x"f4050d74",
   211 => x"53805271",
   212 => x"73259138",
   213 => x"81808051",
   214 => x"c0115170",
   215 => x"fb388112",
   216 => x"5286cf04",
   217 => x"028c050d",
   218 => x"0402f805",
   219 => x"0dec5287",
   220 => x"720c84d8",
   221 => x"5186c72d",
   222 => x"86720c02",
   223 => x"88050d04",
   224 => x"02f8050d",
   225 => x"ec528e72",
   226 => x"0c84d851",
   227 => x"86c72d86",
   228 => x"720c0288",
   229 => x"050d0402",
   230 => x"f8050dec",
   231 => x"5296720c",
   232 => x"84d85186",
   233 => x"c72d8672",
   234 => x"0c028805",
   235 => x"0d0402fc",
   236 => x"050d800b",
   237 => x"bcc00c72",
   238 => x"51b6db2d",
   239 => x"0284050d",
   240 => x"0402fc05",
   241 => x"0d820bbc",
   242 => x"c00c7251",
   243 => x"b6db2d02",
   244 => x"84050d04",
   245 => x"02fc050d",
   246 => x"830bbcc0",
   247 => x"0c7251b6",
   248 => x"db2d0284",
   249 => x"050d0402",
   250 => x"dc050d80",
   251 => x"59a70bec",
   252 => x"0c80e451",
   253 => x"86c72d87",
   254 => x"0bec0c7a",
   255 => x"5280c0f8",
   256 => x"51adf42d",
   257 => x"80c0dc08",
   258 => x"792e80fe",
   259 => x"3880c0fc",
   260 => x"08bcc008",
   261 => x"f00c70f8",
   262 => x"0c79ff12",
   263 => x"56585573",
   264 => x"792e8b38",
   265 => x"81177481",
   266 => x"2a555773",
   267 => x"f738f717",
   268 => x"57815980",
   269 => x"752580d2",
   270 => x"38765273",
   271 => x"5184a82d",
   272 => x"80c1d052",
   273 => x"80c0f851",
   274 => x"b0c12d80",
   275 => x"c0dc0880",
   276 => x"2ea33880",
   277 => x"c1d05880",
   278 => x"56777084",
   279 => x"055908e8",
   280 => x"0cfc1555",
   281 => x"80752595",
   282 => x"38841656",
   283 => x"83ff7625",
   284 => x"e83888fd",
   285 => x"0480c0dc",
   286 => x"0859898a",
   287 => x"0480c0f8",
   288 => x"51b0912d",
   289 => x"81145488",
   290 => x"b304860b",
   291 => x"ec0c7880",
   292 => x"2e9238bc",
   293 => x"c45191bf",
   294 => x"2d8fb72d",
   295 => x"805186e9",
   296 => x"2d89aa04",
   297 => x"beac5191",
   298 => x"bf2d7880",
   299 => x"c0dc0c02",
   300 => x"a4050d04",
   301 => x"02f0050d",
   302 => x"850bec0c",
   303 => x"8ee92d8b",
   304 => x"a12d81f9",
   305 => x"2d83528e",
   306 => x"cc2d8151",
   307 => x"858d2dff",
   308 => x"12527180",
   309 => x"25f138ba",
   310 => x"f05186a0",
   311 => x"2da4b72d",
   312 => x"80c0dc08",
   313 => x"802e81a2",
   314 => x"3887e751",
   315 => x"b6fe2dbc",
   316 => x"c45191bf",
   317 => x"2d8fa42d",
   318 => x"8bad2d91",
   319 => x"d22dbd94",
   320 => x"0b80f52d",
   321 => x"bda00b80",
   322 => x"f52d718a",
   323 => x"2b71832b",
   324 => x"07bdac0b",
   325 => x"80f52d70",
   326 => x"862b7207",
   327 => x"bf980870",
   328 => x"81065354",
   329 => x"52535555",
   330 => x"5271802e",
   331 => x"85387281",
   332 => x"07537381",
   333 => x"2a708106",
   334 => x"51527180",
   335 => x"2e853872",
   336 => x"82075373",
   337 => x"822a7081",
   338 => x"06515271",
   339 => x"802e8538",
   340 => x"72840753",
   341 => x"73832a70",
   342 => x"81065152",
   343 => x"71802e85",
   344 => x"3872a007",
   345 => x"5373842a",
   346 => x"70810651",
   347 => x"5271802e",
   348 => x"86387284",
   349 => x"80075372",
   350 => x"fc0c8652",
   351 => x"80c0dc08",
   352 => x"83388452",
   353 => x"71ec0c89",
   354 => x"f804800b",
   355 => x"80c0dc0c",
   356 => x"0290050d",
   357 => x"0471980c",
   358 => x"04ffb008",
   359 => x"80c0dc0c",
   360 => x"04810bff",
   361 => x"b00c0480",
   362 => x"0bffb00c",
   363 => x"0402f405",
   364 => x"0d80c184",
   365 => x"518db62d",
   366 => x"ff0b80c0",
   367 => x"dc082581",
   368 => x"803880c0",
   369 => x"dc0881f0",
   370 => x"2e098106",
   371 => x"8938810b",
   372 => x"bf900c8c",
   373 => x"c10480c0",
   374 => x"dc0881e0",
   375 => x"2e098106",
   376 => x"8938810b",
   377 => x"bf940c8c",
   378 => x"c10480c0",
   379 => x"dc0852bf",
   380 => x"9408802e",
   381 => x"893880c0",
   382 => x"dc088180",
   383 => x"05527184",
   384 => x"2c728f06",
   385 => x"5353bf90",
   386 => x"08802e99",
   387 => x"38728429",
   388 => x"bed00572",
   389 => x"1381712b",
   390 => x"70097308",
   391 => x"06730c51",
   392 => x"53538cb7",
   393 => x"04728429",
   394 => x"bed00572",
   395 => x"1383712b",
   396 => x"72080772",
   397 => x"0c535380",
   398 => x"0bbf940c",
   399 => x"800bbf90",
   400 => x"0c800b80",
   401 => x"c0dc0c02",
   402 => x"8c050d04",
   403 => x"02f8050d",
   404 => x"bed0528f",
   405 => x"51807270",
   406 => x"8405540c",
   407 => x"ff115170",
   408 => x"8025f238",
   409 => x"0288050d",
   410 => x"0402f005",
   411 => x"0d75518b",
   412 => x"a72d7082",
   413 => x"2cfc06be",
   414 => x"d0117210",
   415 => x"9e067108",
   416 => x"70722a70",
   417 => x"83068274",
   418 => x"2b700974",
   419 => x"06760c54",
   420 => x"51565753",
   421 => x"51538ba1",
   422 => x"2d7180c0",
   423 => x"dc0c0290",
   424 => x"050d0402",
   425 => x"fc050d72",
   426 => x"5180710c",
   427 => x"800b8412",
   428 => x"0c028405",
   429 => x"0d0402f0",
   430 => x"050d7570",
   431 => x"08841208",
   432 => x"535353ff",
   433 => x"5471712e",
   434 => x"a8388ba7",
   435 => x"2d841308",
   436 => x"70842914",
   437 => x"88117008",
   438 => x"7081ff06",
   439 => x"84180881",
   440 => x"11870684",
   441 => x"1a0c5351",
   442 => x"55515151",
   443 => x"8ba12d71",
   444 => x"547380c0",
   445 => x"dc0c0290",
   446 => x"050d0402",
   447 => x"f4050d8b",
   448 => x"a72de008",
   449 => x"708b2a70",
   450 => x"81065152",
   451 => x"5370802e",
   452 => x"a13880c1",
   453 => x"84087084",
   454 => x"2980c18c",
   455 => x"057481ff",
   456 => x"06710c51",
   457 => x"5180c184",
   458 => x"08811187",
   459 => x"0680c184",
   460 => x"0c51728c",
   461 => x"2cbf0680",
   462 => x"c1ac0c80",
   463 => x"0b80c1b0",
   464 => x"0c8b992d",
   465 => x"8ba12d02",
   466 => x"8c050d04",
   467 => x"02fc050d",
   468 => x"8ba72d81",
   469 => x"0b80c1b0",
   470 => x"0c8ba12d",
   471 => x"80c1b008",
   472 => x"5170f938",
   473 => x"0284050d",
   474 => x"0402fc05",
   475 => x"0d80c184",
   476 => x"518da32d",
   477 => x"8ccc2d8d",
   478 => x"fb518b95",
   479 => x"2d028405",
   480 => x"0d0402f8",
   481 => x"050d8fcf",
   482 => x"52815186",
   483 => x"c72dff12",
   484 => x"52718025",
   485 => x"f4380288",
   486 => x"050d0480",
   487 => x"c1bc0880",
   488 => x"c0dc0c04",
   489 => x"02fc050d",
   490 => x"810bbf9c",
   491 => x"0c815185",
   492 => x"8d2d0284",
   493 => x"050d0402",
   494 => x"fc050d8f",
   495 => x"c1048bad",
   496 => x"2d80f651",
   497 => x"8ce92d80",
   498 => x"c0dc08f2",
   499 => x"3880da51",
   500 => x"8ce92d80",
   501 => x"c0dc08e6",
   502 => x"3880c0dc",
   503 => x"08bf9c0c",
   504 => x"80c0dc08",
   505 => x"51858d2d",
   506 => x"0284050d",
   507 => x"0402ec05",
   508 => x"0d765480",
   509 => x"52870b88",
   510 => x"1580f52d",
   511 => x"56537472",
   512 => x"248338a0",
   513 => x"53725183",
   514 => x"842d8112",
   515 => x"8b1580f5",
   516 => x"2d545272",
   517 => x"7225de38",
   518 => x"0294050d",
   519 => x"0402f005",
   520 => x"0d80c1bc",
   521 => x"085481f9",
   522 => x"2d800b80",
   523 => x"c1c00c73",
   524 => x"08802e81",
   525 => x"8538820b",
   526 => x"80c0f00c",
   527 => x"80c1c008",
   528 => x"8f0680c0",
   529 => x"ec0c7308",
   530 => x"5271832e",
   531 => x"96387183",
   532 => x"26893871",
   533 => x"812eaf38",
   534 => x"91a30471",
   535 => x"852e9f38",
   536 => x"91a30488",
   537 => x"1480f52d",
   538 => x"841508bb",
   539 => x"88535452",
   540 => x"86a02d71",
   541 => x"84291370",
   542 => x"08525291",
   543 => x"a7047351",
   544 => x"8fed2d91",
   545 => x"a304bf98",
   546 => x"08881508",
   547 => x"2c708106",
   548 => x"51527180",
   549 => x"2e8738bb",
   550 => x"8c5191a0",
   551 => x"04bb9051",
   552 => x"86a02d84",
   553 => x"14085186",
   554 => x"a02d80c1",
   555 => x"c0088105",
   556 => x"80c1c00c",
   557 => x"8c145490",
   558 => x"af040290",
   559 => x"050d0471",
   560 => x"80c1bc0c",
   561 => x"909d2d80",
   562 => x"c1c008ff",
   563 => x"0580c1c4",
   564 => x"0c0402e8",
   565 => x"050d80c1",
   566 => x"bc0880c1",
   567 => x"c8085755",
   568 => x"80f6518c",
   569 => x"e92d80c0",
   570 => x"dc08812a",
   571 => x"70810651",
   572 => x"5271802e",
   573 => x"a03891fc",
   574 => x"048bad2d",
   575 => x"80f6518c",
   576 => x"e92d80c0",
   577 => x"dc08f238",
   578 => x"bf9c0881",
   579 => x"3270bf9c",
   580 => x"0c51858d",
   581 => x"2d80c1ac",
   582 => x"08a00652",
   583 => x"80722596",
   584 => x"388f822d",
   585 => x"8bad2dbf",
   586 => x"9c088132",
   587 => x"70bf9c0c",
   588 => x"70525285",
   589 => x"8d2d800b",
   590 => x"80c1b40c",
   591 => x"800b80c1",
   592 => x"b80cbf9c",
   593 => x"0883ad38",
   594 => x"80da518c",
   595 => x"e92d80c0",
   596 => x"dc08802e",
   597 => x"8c3880c1",
   598 => x"b4088180",
   599 => x"0780c1b4",
   600 => x"0c80d951",
   601 => x"8ce92d80",
   602 => x"c0dc0880",
   603 => x"2e8c3880",
   604 => x"c1b40880",
   605 => x"c00780c1",
   606 => x"b40c8194",
   607 => x"518ce92d",
   608 => x"80c0dc08",
   609 => x"802e8b38",
   610 => x"80c1b408",
   611 => x"900780c1",
   612 => x"b40c8191",
   613 => x"518ce92d",
   614 => x"80c0dc08",
   615 => x"802e8b38",
   616 => x"80c1b408",
   617 => x"a00780c1",
   618 => x"b40c81f5",
   619 => x"518ce92d",
   620 => x"80c0dc08",
   621 => x"802e8b38",
   622 => x"80c1b408",
   623 => x"810780c1",
   624 => x"b40c81f2",
   625 => x"518ce92d",
   626 => x"80c0dc08",
   627 => x"802e8b38",
   628 => x"80c1b408",
   629 => x"820780c1",
   630 => x"b40c81eb",
   631 => x"518ce92d",
   632 => x"80c0dc08",
   633 => x"802e8b38",
   634 => x"80c1b408",
   635 => x"840780c1",
   636 => x"b40c81f4",
   637 => x"518ce92d",
   638 => x"80c0dc08",
   639 => x"802e8b38",
   640 => x"80c1b408",
   641 => x"880780c1",
   642 => x"b40c80d8",
   643 => x"518ce92d",
   644 => x"80c0dc08",
   645 => x"802e8c38",
   646 => x"80c1b808",
   647 => x"81800780",
   648 => x"c1b80c92",
   649 => x"518ce92d",
   650 => x"80c0dc08",
   651 => x"802e8c38",
   652 => x"80c1b808",
   653 => x"80c00780",
   654 => x"c1b80c94",
   655 => x"518ce92d",
   656 => x"80c0dc08",
   657 => x"802e8b38",
   658 => x"80c1b808",
   659 => x"900780c1",
   660 => x"b80c9151",
   661 => x"8ce92d80",
   662 => x"c0dc0880",
   663 => x"2e8b3880",
   664 => x"c1b808a0",
   665 => x"0780c1b8",
   666 => x"0c9d518c",
   667 => x"e92d80c0",
   668 => x"dc08802e",
   669 => x"8b3880c1",
   670 => x"b8088107",
   671 => x"80c1b80c",
   672 => x"9b518ce9",
   673 => x"2d80c0dc",
   674 => x"08802e8b",
   675 => x"3880c1b8",
   676 => x"08820780",
   677 => x"c1b80c9c",
   678 => x"518ce92d",
   679 => x"80c0dc08",
   680 => x"802e8b38",
   681 => x"80c1b808",
   682 => x"840780c1",
   683 => x"b80ca351",
   684 => x"8ce92d80",
   685 => x"c0dc0880",
   686 => x"2e8b3880",
   687 => x"c1b80888",
   688 => x"0780c1b8",
   689 => x"0c96518c",
   690 => x"e92d80c0",
   691 => x"dc08802e",
   692 => x"84388797",
   693 => x"2d9e518c",
   694 => x"e92d80c0",
   695 => x"dc08802e",
   696 => x"84388780",
   697 => x"2d81fd51",
   698 => x"8ce92d81",
   699 => x"fa518ce9",
   700 => x"2d9c9304",
   701 => x"81f5518c",
   702 => x"e92d80c0",
   703 => x"dc08812a",
   704 => x"70810651",
   705 => x"52718e38",
   706 => x"80c1ac08",
   707 => x"90065280",
   708 => x"722580c2",
   709 => x"3880c1ac",
   710 => x"08900652",
   711 => x"80722584",
   712 => x"388f822d",
   713 => x"80c1c408",
   714 => x"5271802e",
   715 => x"8a38ff12",
   716 => x"80c1c40c",
   717 => x"96d60480",
   718 => x"c1c00810",
   719 => x"80c1c008",
   720 => x"05708429",
   721 => x"16515288",
   722 => x"1208802e",
   723 => x"8938ff51",
   724 => x"88120852",
   725 => x"712d81f2",
   726 => x"518ce92d",
   727 => x"80c0dc08",
   728 => x"812a7081",
   729 => x"06515271",
   730 => x"8e3880c1",
   731 => x"ac088806",
   732 => x"52807225",
   733 => x"80c33880",
   734 => x"c1ac0888",
   735 => x"06528072",
   736 => x"2584388f",
   737 => x"822d80c1",
   738 => x"c008ff11",
   739 => x"80c1c408",
   740 => x"56535373",
   741 => x"72258a38",
   742 => x"811480c1",
   743 => x"c40c97b9",
   744 => x"04721013",
   745 => x"70842916",
   746 => x"51528812",
   747 => x"08802e89",
   748 => x"38fe5188",
   749 => x"12085271",
   750 => x"2d81fd51",
   751 => x"8ce92d80",
   752 => x"c0dc0881",
   753 => x"2a708106",
   754 => x"51527180",
   755 => x"2eb13880",
   756 => x"c1c40880",
   757 => x"2e8a3880",
   758 => x"0b80c1c4",
   759 => x"0c97ff04",
   760 => x"80c1c008",
   761 => x"1080c1c0",
   762 => x"08057084",
   763 => x"29165152",
   764 => x"88120880",
   765 => x"2e8938fd",
   766 => x"51881208",
   767 => x"52712d81",
   768 => x"fa518ce9",
   769 => x"2d80c0dc",
   770 => x"08812a70",
   771 => x"81065152",
   772 => x"71802eb1",
   773 => x"3880c1c0",
   774 => x"08ff1154",
   775 => x"5280c1c4",
   776 => x"08732589",
   777 => x"387280c1",
   778 => x"c40c98c5",
   779 => x"04711012",
   780 => x"70842916",
   781 => x"51528812",
   782 => x"08802e89",
   783 => x"38fc5188",
   784 => x"12085271",
   785 => x"2d80c1c4",
   786 => x"08705354",
   787 => x"73802e8a",
   788 => x"388c15ff",
   789 => x"15555598",
   790 => x"cc04820b",
   791 => x"80c0f00c",
   792 => x"718f0680",
   793 => x"c0ec0c81",
   794 => x"eb518ce9",
   795 => x"2d80c0dc",
   796 => x"08812a70",
   797 => x"81065152",
   798 => x"71802ead",
   799 => x"38740885",
   800 => x"2e098106",
   801 => x"a4388815",
   802 => x"80f52dff",
   803 => x"05527188",
   804 => x"1681b72d",
   805 => x"71982b52",
   806 => x"71802588",
   807 => x"38800b88",
   808 => x"1681b72d",
   809 => x"74518fed",
   810 => x"2d81f451",
   811 => x"8ce92d80",
   812 => x"c0dc0881",
   813 => x"2a708106",
   814 => x"51527180",
   815 => x"2eb33874",
   816 => x"08852e09",
   817 => x"8106aa38",
   818 => x"881580f5",
   819 => x"2d810552",
   820 => x"71881681",
   821 => x"b72d7181",
   822 => x"ff068b16",
   823 => x"80f52d54",
   824 => x"52727227",
   825 => x"87387288",
   826 => x"1681b72d",
   827 => x"74518fed",
   828 => x"2d80da51",
   829 => x"8ce92d80",
   830 => x"c0dc0881",
   831 => x"2a708106",
   832 => x"5152718e",
   833 => x"3880c1ac",
   834 => x"08810652",
   835 => x"80722581",
   836 => x"ba3880c1",
   837 => x"bc0880c1",
   838 => x"ac088106",
   839 => x"53538072",
   840 => x"2584388f",
   841 => x"822d80c1",
   842 => x"c4085473",
   843 => x"802e8a38",
   844 => x"8c13ff15",
   845 => x"55539aab",
   846 => x"04720852",
   847 => x"71822ea6",
   848 => x"38718226",
   849 => x"89387181",
   850 => x"2eaa389b",
   851 => x"cb047183",
   852 => x"2eb23871",
   853 => x"842e0981",
   854 => x"0680f038",
   855 => x"88130851",
   856 => x"91bf2d9b",
   857 => x"cb0480c1",
   858 => x"c4085188",
   859 => x"13085271",
   860 => x"2d9bcb04",
   861 => x"810b8814",
   862 => x"082bbf98",
   863 => x"0832bf98",
   864 => x"0c9b9f04",
   865 => x"881380f5",
   866 => x"2d81058b",
   867 => x"1480f52d",
   868 => x"53547174",
   869 => x"24833880",
   870 => x"54738814",
   871 => x"81b72d90",
   872 => x"9d2d9bcb",
   873 => x"04750880",
   874 => x"2ea43875",
   875 => x"08518ce9",
   876 => x"2d80c0dc",
   877 => x"08810652",
   878 => x"71802e8c",
   879 => x"3880c1c4",
   880 => x"08518416",
   881 => x"0852712d",
   882 => x"88165675",
   883 => x"d8388054",
   884 => x"800b80c0",
   885 => x"f00c738f",
   886 => x"0680c0ec",
   887 => x"0ca05273",
   888 => x"80c1c408",
   889 => x"2e098106",
   890 => x"993880c1",
   891 => x"c008ff05",
   892 => x"74327009",
   893 => x"81057072",
   894 => x"079f2a91",
   895 => x"71315151",
   896 => x"53537151",
   897 => x"83842d81",
   898 => x"14548e74",
   899 => x"25c238bf",
   900 => x"9c085271",
   901 => x"80c0dc0c",
   902 => x"0298050d",
   903 => x"0402f405",
   904 => x"0dd45281",
   905 => x"ff720c71",
   906 => x"085381ff",
   907 => x"720c7288",
   908 => x"2b83fe80",
   909 => x"06720870",
   910 => x"81ff0651",
   911 => x"525381ff",
   912 => x"720c7271",
   913 => x"07882b72",
   914 => x"087081ff",
   915 => x"06515253",
   916 => x"81ff720c",
   917 => x"72710788",
   918 => x"2b720870",
   919 => x"81ff0672",
   920 => x"0780c0dc",
   921 => x"0c525302",
   922 => x"8c050d04",
   923 => x"02f4050d",
   924 => x"74767181",
   925 => x"ff06d40c",
   926 => x"535380c1",
   927 => x"cc088538",
   928 => x"71892b52",
   929 => x"71982ad4",
   930 => x"0c71902a",
   931 => x"7081ff06",
   932 => x"d40c5171",
   933 => x"882a7081",
   934 => x"ff06d40c",
   935 => x"517181ff",
   936 => x"06d40c72",
   937 => x"902a7081",
   938 => x"ff06d40c",
   939 => x"51d40870",
   940 => x"81ff0651",
   941 => x"5182b8bf",
   942 => x"527081ff",
   943 => x"2e098106",
   944 => x"943881ff",
   945 => x"0bd40cd4",
   946 => x"087081ff",
   947 => x"06ff1454",
   948 => x"515171e5",
   949 => x"387080c0",
   950 => x"dc0c028c",
   951 => x"050d0402",
   952 => x"fc050d81",
   953 => x"c75181ff",
   954 => x"0bd40cff",
   955 => x"11517080",
   956 => x"25f43802",
   957 => x"84050d04",
   958 => x"02f4050d",
   959 => x"81ff0bd4",
   960 => x"0c935380",
   961 => x"5287fc80",
   962 => x"c1519cec",
   963 => x"2d80c0dc",
   964 => x"088b3881",
   965 => x"ff0bd40c",
   966 => x"81539ea6",
   967 => x"049ddf2d",
   968 => x"ff135372",
   969 => x"de387280",
   970 => x"c0dc0c02",
   971 => x"8c050d04",
   972 => x"02ec050d",
   973 => x"810b80c1",
   974 => x"cc0c8454",
   975 => x"d008708f",
   976 => x"2a708106",
   977 => x"51515372",
   978 => x"f33872d0",
   979 => x"0c9ddf2d",
   980 => x"bb945186",
   981 => x"a02dd008",
   982 => x"708f2a70",
   983 => x"81065151",
   984 => x"5372f338",
   985 => x"810bd00c",
   986 => x"b1538052",
   987 => x"84d480c0",
   988 => x"519cec2d",
   989 => x"80c0dc08",
   990 => x"812e9338",
   991 => x"72822ebf",
   992 => x"38ff1353",
   993 => x"72e438ff",
   994 => x"145473ff",
   995 => x"af389ddf",
   996 => x"2d83aa52",
   997 => x"849c80c8",
   998 => x"519cec2d",
   999 => x"80c0dc08",
  1000 => x"812e0981",
  1001 => x"0693389c",
  1002 => x"9d2d80c0",
  1003 => x"dc0883ff",
  1004 => x"ff065372",
  1005 => x"83aa2e9d",
  1006 => x"389df82d",
  1007 => x"9fd004bb",
  1008 => x"a05186a0",
  1009 => x"2d8053a1",
  1010 => x"a504bbb8",
  1011 => x"5186a02d",
  1012 => x"8054a0f6",
  1013 => x"0481ff0b",
  1014 => x"d40cb154",
  1015 => x"9ddf2d8f",
  1016 => x"cf538052",
  1017 => x"87fc80f7",
  1018 => x"519cec2d",
  1019 => x"80c0dc08",
  1020 => x"5580c0dc",
  1021 => x"08812e09",
  1022 => x"81069c38",
  1023 => x"81ff0bd4",
  1024 => x"0c820a52",
  1025 => x"849c80e9",
  1026 => x"519cec2d",
  1027 => x"80c0dc08",
  1028 => x"802e8d38",
  1029 => x"9ddf2dff",
  1030 => x"135372c6",
  1031 => x"38a0e904",
  1032 => x"81ff0bd4",
  1033 => x"0c80c0dc",
  1034 => x"085287fc",
  1035 => x"80fa519c",
  1036 => x"ec2d80c0",
  1037 => x"dc08b238",
  1038 => x"81ff0bd4",
  1039 => x"0cd40853",
  1040 => x"81ff0bd4",
  1041 => x"0c81ff0b",
  1042 => x"d40c81ff",
  1043 => x"0bd40c81",
  1044 => x"ff0bd40c",
  1045 => x"72862a70",
  1046 => x"81067656",
  1047 => x"51537296",
  1048 => x"3880c0dc",
  1049 => x"0854a0f6",
  1050 => x"0473822e",
  1051 => x"fedc38ff",
  1052 => x"145473fe",
  1053 => x"e7387380",
  1054 => x"c1cc0c73",
  1055 => x"8b388152",
  1056 => x"87fc80d0",
  1057 => x"519cec2d",
  1058 => x"81ff0bd4",
  1059 => x"0cd00870",
  1060 => x"8f2a7081",
  1061 => x"06515153",
  1062 => x"72f33872",
  1063 => x"d00c81ff",
  1064 => x"0bd40c81",
  1065 => x"537280c0",
  1066 => x"dc0c0294",
  1067 => x"050d0402",
  1068 => x"e8050d78",
  1069 => x"55805681",
  1070 => x"ff0bd40c",
  1071 => x"d008708f",
  1072 => x"2a708106",
  1073 => x"51515372",
  1074 => x"f3388281",
  1075 => x"0bd00c81",
  1076 => x"ff0bd40c",
  1077 => x"775287fc",
  1078 => x"80d1519c",
  1079 => x"ec2d80db",
  1080 => x"c6df5480",
  1081 => x"c0dc0880",
  1082 => x"2e8a38bb",
  1083 => x"d85186a0",
  1084 => x"2da2c804",
  1085 => x"81ff0bd4",
  1086 => x"0cd40870",
  1087 => x"81ff0651",
  1088 => x"537281fe",
  1089 => x"2e098106",
  1090 => x"9e3880ff",
  1091 => x"539c9d2d",
  1092 => x"80c0dc08",
  1093 => x"75708405",
  1094 => x"570cff13",
  1095 => x"53728025",
  1096 => x"ec388156",
  1097 => x"a2ad04ff",
  1098 => x"145473c8",
  1099 => x"3881ff0b",
  1100 => x"d40c81ff",
  1101 => x"0bd40cd0",
  1102 => x"08708f2a",
  1103 => x"70810651",
  1104 => x"515372f3",
  1105 => x"3872d00c",
  1106 => x"7580c0dc",
  1107 => x"0c029805",
  1108 => x"0d0402e8",
  1109 => x"050d7779",
  1110 => x"7b585555",
  1111 => x"80537276",
  1112 => x"25a33874",
  1113 => x"70810556",
  1114 => x"80f52d74",
  1115 => x"70810556",
  1116 => x"80f52d52",
  1117 => x"5271712e",
  1118 => x"86388151",
  1119 => x"a3870481",
  1120 => x"1353a2de",
  1121 => x"04805170",
  1122 => x"80c0dc0c",
  1123 => x"0298050d",
  1124 => x"0402ec05",
  1125 => x"0d765574",
  1126 => x"802e80c2",
  1127 => x"389a1580",
  1128 => x"e02d51b1",
  1129 => x"9b2d80c0",
  1130 => x"dc0880c0",
  1131 => x"dc0880c8",
  1132 => x"800c80c0",
  1133 => x"dc085454",
  1134 => x"80c7dc08",
  1135 => x"802e9a38",
  1136 => x"941580e0",
  1137 => x"2d51b19b",
  1138 => x"2d80c0dc",
  1139 => x"08902b83",
  1140 => x"fff00a06",
  1141 => x"70750751",
  1142 => x"537280c8",
  1143 => x"800c80c8",
  1144 => x"80085372",
  1145 => x"802e9d38",
  1146 => x"80c7d408",
  1147 => x"fe147129",
  1148 => x"80c7e808",
  1149 => x"0580c884",
  1150 => x"0c70842b",
  1151 => x"80c7e00c",
  1152 => x"54a4b204",
  1153 => x"80c7ec08",
  1154 => x"80c8800c",
  1155 => x"80c7f008",
  1156 => x"80c8840c",
  1157 => x"80c7dc08",
  1158 => x"802e8b38",
  1159 => x"80c7d408",
  1160 => x"842b53a4",
  1161 => x"ad0480c7",
  1162 => x"f408842b",
  1163 => x"537280c7",
  1164 => x"e00c0294",
  1165 => x"050d0402",
  1166 => x"d8050d80",
  1167 => x"0b80c7dc",
  1168 => x"0c84549e",
  1169 => x"b02d80c0",
  1170 => x"dc08802e",
  1171 => x"973880c1",
  1172 => x"d0528051",
  1173 => x"a1af2d80",
  1174 => x"c0dc0880",
  1175 => x"2e8638fe",
  1176 => x"54a4ec04",
  1177 => x"ff145473",
  1178 => x"8024d838",
  1179 => x"738c38bb",
  1180 => x"e85186a0",
  1181 => x"2d7355aa",
  1182 => x"b9048056",
  1183 => x"810b80c8",
  1184 => x"880c8853",
  1185 => x"bbfc5280",
  1186 => x"c28651a2",
  1187 => x"d22d80c0",
  1188 => x"dc08762e",
  1189 => x"09810689",
  1190 => x"3880c0dc",
  1191 => x"0880c888",
  1192 => x"0c8853bc",
  1193 => x"885280c2",
  1194 => x"a251a2d2",
  1195 => x"2d80c0dc",
  1196 => x"08893880",
  1197 => x"c0dc0880",
  1198 => x"c8880c80",
  1199 => x"c8880880",
  1200 => x"2e818038",
  1201 => x"80c5960b",
  1202 => x"80f52d80",
  1203 => x"c5970b80",
  1204 => x"f52d7198",
  1205 => x"2b71902b",
  1206 => x"0780c598",
  1207 => x"0b80f52d",
  1208 => x"70882b72",
  1209 => x"0780c599",
  1210 => x"0b80f52d",
  1211 => x"710780c5",
  1212 => x"ce0b80f5",
  1213 => x"2d80c5cf",
  1214 => x"0b80f52d",
  1215 => x"71882b07",
  1216 => x"535f5452",
  1217 => x"5a565755",
  1218 => x"7381abaa",
  1219 => x"2e098106",
  1220 => x"8e387551",
  1221 => x"b0ea2d80",
  1222 => x"c0dc0856",
  1223 => x"a6ac0473",
  1224 => x"82d4d52e",
  1225 => x"8738bc94",
  1226 => x"51a6f504",
  1227 => x"80c1d052",
  1228 => x"7551a1af",
  1229 => x"2d80c0dc",
  1230 => x"085580c0",
  1231 => x"dc08802e",
  1232 => x"83f73888",
  1233 => x"53bc8852",
  1234 => x"80c2a251",
  1235 => x"a2d22d80",
  1236 => x"c0dc088a",
  1237 => x"38810b80",
  1238 => x"c7dc0ca6",
  1239 => x"fb048853",
  1240 => x"bbfc5280",
  1241 => x"c28651a2",
  1242 => x"d22d80c0",
  1243 => x"dc08802e",
  1244 => x"8a38bca8",
  1245 => x"5186a02d",
  1246 => x"a7da0480",
  1247 => x"c5ce0b80",
  1248 => x"f52d5473",
  1249 => x"80d52e09",
  1250 => x"810680ce",
  1251 => x"3880c5cf",
  1252 => x"0b80f52d",
  1253 => x"547381aa",
  1254 => x"2e098106",
  1255 => x"bd38800b",
  1256 => x"80c1d00b",
  1257 => x"80f52d56",
  1258 => x"547481e9",
  1259 => x"2e833881",
  1260 => x"547481eb",
  1261 => x"2e8c3880",
  1262 => x"5573752e",
  1263 => x"09810682",
  1264 => x"f83880c1",
  1265 => x"db0b80f5",
  1266 => x"2d55748e",
  1267 => x"3880c1dc",
  1268 => x"0b80f52d",
  1269 => x"5473822e",
  1270 => x"86388055",
  1271 => x"aab90480",
  1272 => x"c1dd0b80",
  1273 => x"f52d7080",
  1274 => x"c7d40cff",
  1275 => x"0580c7d8",
  1276 => x"0c80c1de",
  1277 => x"0b80f52d",
  1278 => x"80c1df0b",
  1279 => x"80f52d58",
  1280 => x"76057782",
  1281 => x"80290570",
  1282 => x"80c7e40c",
  1283 => x"80c1e00b",
  1284 => x"80f52d70",
  1285 => x"80c7f80c",
  1286 => x"80c7dc08",
  1287 => x"59575876",
  1288 => x"802e81b6",
  1289 => x"388853bc",
  1290 => x"885280c2",
  1291 => x"a251a2d2",
  1292 => x"2d80c0dc",
  1293 => x"08828238",
  1294 => x"80c7d408",
  1295 => x"70842b80",
  1296 => x"c7e00c70",
  1297 => x"80c7f40c",
  1298 => x"80c1f50b",
  1299 => x"80f52d80",
  1300 => x"c1f40b80",
  1301 => x"f52d7182",
  1302 => x"80290580",
  1303 => x"c1f60b80",
  1304 => x"f52d7084",
  1305 => x"80802912",
  1306 => x"80c1f70b",
  1307 => x"80f52d70",
  1308 => x"81800a29",
  1309 => x"127080c7",
  1310 => x"fc0c80c7",
  1311 => x"f8087129",
  1312 => x"80c7e408",
  1313 => x"057080c7",
  1314 => x"e80c80c1",
  1315 => x"fd0b80f5",
  1316 => x"2d80c1fc",
  1317 => x"0b80f52d",
  1318 => x"71828029",
  1319 => x"0580c1fe",
  1320 => x"0b80f52d",
  1321 => x"70848080",
  1322 => x"291280c1",
  1323 => x"ff0b80f5",
  1324 => x"2d70982b",
  1325 => x"81f00a06",
  1326 => x"72057080",
  1327 => x"c7ec0cfe",
  1328 => x"117e2977",
  1329 => x"0580c7f0",
  1330 => x"0c525952",
  1331 => x"43545e51",
  1332 => x"5259525d",
  1333 => x"575957aa",
  1334 => x"b20480c1",
  1335 => x"e20b80f5",
  1336 => x"2d80c1e1",
  1337 => x"0b80f52d",
  1338 => x"71828029",
  1339 => x"057080c7",
  1340 => x"e00c70a0",
  1341 => x"2983ff05",
  1342 => x"70892a70",
  1343 => x"80c7f40c",
  1344 => x"80c1e70b",
  1345 => x"80f52d80",
  1346 => x"c1e60b80",
  1347 => x"f52d7182",
  1348 => x"80290570",
  1349 => x"80c7fc0c",
  1350 => x"7b71291e",
  1351 => x"7080c7f0",
  1352 => x"0c7d80c7",
  1353 => x"ec0c7305",
  1354 => x"80c7e80c",
  1355 => x"555e5151",
  1356 => x"55558051",
  1357 => x"a3912d81",
  1358 => x"557480c0",
  1359 => x"dc0c02a8",
  1360 => x"050d0402",
  1361 => x"ec050d76",
  1362 => x"70872c71",
  1363 => x"80ff0655",
  1364 => x"565480c7",
  1365 => x"dc088a38",
  1366 => x"73882c74",
  1367 => x"81ff0654",
  1368 => x"5580c1d0",
  1369 => x"5280c7e4",
  1370 => x"081551a1",
  1371 => x"af2d80c0",
  1372 => x"dc085480",
  1373 => x"c0dc0880",
  1374 => x"2eb83880",
  1375 => x"c7dc0880",
  1376 => x"2e9a3872",
  1377 => x"842980c1",
  1378 => x"d0057008",
  1379 => x"5253b0ea",
  1380 => x"2d80c0dc",
  1381 => x"08f00a06",
  1382 => x"53abb004",
  1383 => x"721080c1",
  1384 => x"d0057080",
  1385 => x"e02d5253",
  1386 => x"b19b2d80",
  1387 => x"c0dc0853",
  1388 => x"72547380",
  1389 => x"c0dc0c02",
  1390 => x"94050d04",
  1391 => x"02e0050d",
  1392 => x"7970842c",
  1393 => x"80c88408",
  1394 => x"05718f06",
  1395 => x"52555372",
  1396 => x"8a3880c1",
  1397 => x"d0527351",
  1398 => x"a1af2d72",
  1399 => x"a02980c1",
  1400 => x"d0055480",
  1401 => x"7480f52d",
  1402 => x"56537473",
  1403 => x"2e833881",
  1404 => x"537481e5",
  1405 => x"2e81f138",
  1406 => x"81707406",
  1407 => x"54587280",
  1408 => x"2e81e538",
  1409 => x"8b1480f5",
  1410 => x"2d70832a",
  1411 => x"79065856",
  1412 => x"769938bf",
  1413 => x"a0085372",
  1414 => x"89387280",
  1415 => x"c5d00b81",
  1416 => x"b72d76bf",
  1417 => x"a00c7353",
  1418 => x"adea0475",
  1419 => x"8f2e0981",
  1420 => x"0681b538",
  1421 => x"749f068d",
  1422 => x"2980c5c3",
  1423 => x"11515381",
  1424 => x"1480f52d",
  1425 => x"73708105",
  1426 => x"5581b72d",
  1427 => x"831480f5",
  1428 => x"2d737081",
  1429 => x"055581b7",
  1430 => x"2d851480",
  1431 => x"f52d7370",
  1432 => x"81055581",
  1433 => x"b72d8714",
  1434 => x"80f52d73",
  1435 => x"70810555",
  1436 => x"81b72d89",
  1437 => x"1480f52d",
  1438 => x"73708105",
  1439 => x"5581b72d",
  1440 => x"8e1480f5",
  1441 => x"2d737081",
  1442 => x"055581b7",
  1443 => x"2d901480",
  1444 => x"f52d7370",
  1445 => x"81055581",
  1446 => x"b72d9214",
  1447 => x"80f52d73",
  1448 => x"70810555",
  1449 => x"81b72d94",
  1450 => x"1480f52d",
  1451 => x"73708105",
  1452 => x"5581b72d",
  1453 => x"961480f5",
  1454 => x"2d737081",
  1455 => x"055581b7",
  1456 => x"2d981480",
  1457 => x"f52d7370",
  1458 => x"81055581",
  1459 => x"b72d9c14",
  1460 => x"80f52d73",
  1461 => x"70810555",
  1462 => x"81b72d9e",
  1463 => x"1480f52d",
  1464 => x"7381b72d",
  1465 => x"77bfa00c",
  1466 => x"80537280",
  1467 => x"c0dc0c02",
  1468 => x"a0050d04",
  1469 => x"02cc050d",
  1470 => x"7e605e5a",
  1471 => x"800b80c8",
  1472 => x"800880c8",
  1473 => x"8408595c",
  1474 => x"56805880",
  1475 => x"c7e00878",
  1476 => x"2e81b838",
  1477 => x"778f06a0",
  1478 => x"17575473",
  1479 => x"913880c1",
  1480 => x"d0527651",
  1481 => x"811757a1",
  1482 => x"af2d80c1",
  1483 => x"d0568076",
  1484 => x"80f52d56",
  1485 => x"5474742e",
  1486 => x"83388154",
  1487 => x"7481e52e",
  1488 => x"80fd3881",
  1489 => x"70750655",
  1490 => x"5c73802e",
  1491 => x"80f1388b",
  1492 => x"1680f52d",
  1493 => x"98065978",
  1494 => x"80e5388b",
  1495 => x"537c5275",
  1496 => x"51a2d22d",
  1497 => x"80c0dc08",
  1498 => x"80d5389c",
  1499 => x"160851b0",
  1500 => x"ea2d80c0",
  1501 => x"dc08841b",
  1502 => x"0c9a1680",
  1503 => x"e02d51b1",
  1504 => x"9b2d80c0",
  1505 => x"dc0880c0",
  1506 => x"dc08881c",
  1507 => x"0c80c0dc",
  1508 => x"08555580",
  1509 => x"c7dc0880",
  1510 => x"2e993894",
  1511 => x"1680e02d",
  1512 => x"51b19b2d",
  1513 => x"80c0dc08",
  1514 => x"902b83ff",
  1515 => x"f00a0670",
  1516 => x"16515473",
  1517 => x"881b0c78",
  1518 => x"7a0c7b54",
  1519 => x"b0870481",
  1520 => x"185880c7",
  1521 => x"e0087826",
  1522 => x"feca3880",
  1523 => x"c7dc0880",
  1524 => x"2eb3387a",
  1525 => x"51aac32d",
  1526 => x"80c0dc08",
  1527 => x"80c0dc08",
  1528 => x"80ffffff",
  1529 => x"f806555b",
  1530 => x"7380ffff",
  1531 => x"fff82e95",
  1532 => x"3880c0dc",
  1533 => x"08fe0580",
  1534 => x"c7d40829",
  1535 => x"80c7e808",
  1536 => x"0557ae89",
  1537 => x"04805473",
  1538 => x"80c0dc0c",
  1539 => x"02b4050d",
  1540 => x"0402f405",
  1541 => x"0d747008",
  1542 => x"8105710c",
  1543 => x"700880c7",
  1544 => x"d8080653",
  1545 => x"53718f38",
  1546 => x"88130851",
  1547 => x"aac32d80",
  1548 => x"c0dc0888",
  1549 => x"140c810b",
  1550 => x"80c0dc0c",
  1551 => x"028c050d",
  1552 => x"0402f005",
  1553 => x"0d758811",
  1554 => x"08fe0580",
  1555 => x"c7d40829",
  1556 => x"80c7e808",
  1557 => x"11720880",
  1558 => x"c7d80806",
  1559 => x"05795553",
  1560 => x"5454a1af",
  1561 => x"2d029005",
  1562 => x"0d0402f4",
  1563 => x"050d7470",
  1564 => x"882a83fe",
  1565 => x"80067072",
  1566 => x"982a0772",
  1567 => x"882b87fc",
  1568 => x"80800673",
  1569 => x"982b81f0",
  1570 => x"0a067173",
  1571 => x"070780c0",
  1572 => x"dc0c5651",
  1573 => x"5351028c",
  1574 => x"050d0402",
  1575 => x"f8050d02",
  1576 => x"8e0580f5",
  1577 => x"2d74882b",
  1578 => x"077083ff",
  1579 => x"ff0680c0",
  1580 => x"dc0c5102",
  1581 => x"88050d04",
  1582 => x"02f4050d",
  1583 => x"74767853",
  1584 => x"54528071",
  1585 => x"25973872",
  1586 => x"70810554",
  1587 => x"80f52d72",
  1588 => x"70810554",
  1589 => x"81b72dff",
  1590 => x"115170eb",
  1591 => x"38807281",
  1592 => x"b72d028c",
  1593 => x"050d0402",
  1594 => x"e8050d77",
  1595 => x"56807056",
  1596 => x"54737624",
  1597 => x"b63880c7",
  1598 => x"e008742e",
  1599 => x"ae387351",
  1600 => x"abbc2d80",
  1601 => x"c0dc0880",
  1602 => x"c0dc0809",
  1603 => x"81057080",
  1604 => x"c0dc0807",
  1605 => x"9f2a7705",
  1606 => x"81175757",
  1607 => x"53537476",
  1608 => x"24893880",
  1609 => x"c7e00874",
  1610 => x"26d43872",
  1611 => x"80c0dc0c",
  1612 => x"0298050d",
  1613 => x"0402f005",
  1614 => x"0d80c0d8",
  1615 => x"081651b1",
  1616 => x"e72d80c0",
  1617 => x"dc08802e",
  1618 => x"9f388b53",
  1619 => x"80c0dc08",
  1620 => x"5280c5d0",
  1621 => x"51b1b82d",
  1622 => x"80c88c08",
  1623 => x"5473802e",
  1624 => x"873880c5",
  1625 => x"d051732d",
  1626 => x"0290050d",
  1627 => x"0402dc05",
  1628 => x"0d80705a",
  1629 => x"557480c0",
  1630 => x"d80825b4",
  1631 => x"3880c7e0",
  1632 => x"08752eac",
  1633 => x"387851ab",
  1634 => x"bc2d80c0",
  1635 => x"dc080981",
  1636 => x"057080c0",
  1637 => x"dc08079f",
  1638 => x"2a760581",
  1639 => x"1b5b5654",
  1640 => x"7480c0d8",
  1641 => x"08258938",
  1642 => x"80c7e008",
  1643 => x"7926d638",
  1644 => x"80557880",
  1645 => x"c7e00827",
  1646 => x"81d93878",
  1647 => x"51abbc2d",
  1648 => x"80c0dc08",
  1649 => x"802e81ab",
  1650 => x"3880c0dc",
  1651 => x"088b0580",
  1652 => x"f52d7084",
  1653 => x"2a708106",
  1654 => x"77107884",
  1655 => x"2b80c5d0",
  1656 => x"0b80f52d",
  1657 => x"5c5c5351",
  1658 => x"55567380",
  1659 => x"2e80ca38",
  1660 => x"7416822b",
  1661 => x"b5b70bbf",
  1662 => x"ac120c54",
  1663 => x"77753110",
  1664 => x"80c89011",
  1665 => x"55569074",
  1666 => x"70810556",
  1667 => x"81b72da0",
  1668 => x"7481b72d",
  1669 => x"7681ff06",
  1670 => x"81165854",
  1671 => x"73802e8a",
  1672 => x"389c5380",
  1673 => x"c5d052b4",
  1674 => x"b1048b53",
  1675 => x"80c0dc08",
  1676 => x"5280c892",
  1677 => x"1651b4eb",
  1678 => x"04741682",
  1679 => x"2bb2b50b",
  1680 => x"bfac120c",
  1681 => x"547681ff",
  1682 => x"06811658",
  1683 => x"5473802e",
  1684 => x"8a389c53",
  1685 => x"80c5d052",
  1686 => x"b4e2048b",
  1687 => x"5380c0dc",
  1688 => x"08527775",
  1689 => x"311080c8",
  1690 => x"90055176",
  1691 => x"55b1b82d",
  1692 => x"b5880474",
  1693 => x"90297531",
  1694 => x"701080c8",
  1695 => x"90055154",
  1696 => x"80c0dc08",
  1697 => x"7481b72d",
  1698 => x"81195974",
  1699 => x"8b24a338",
  1700 => x"b3b20474",
  1701 => x"90297531",
  1702 => x"701080c8",
  1703 => x"90058c77",
  1704 => x"31575154",
  1705 => x"807481b7",
  1706 => x"2d9e14ff",
  1707 => x"16565474",
  1708 => x"f33802a4",
  1709 => x"050d0402",
  1710 => x"fc050d80",
  1711 => x"c0d80813",
  1712 => x"51b1e72d",
  1713 => x"80c0dc08",
  1714 => x"802e8938",
  1715 => x"80c0dc08",
  1716 => x"51a3912d",
  1717 => x"800b80c0",
  1718 => x"d80cb2ed",
  1719 => x"2d909d2d",
  1720 => x"0284050d",
  1721 => x"0402fc05",
  1722 => x"0d725170",
  1723 => x"fd2eb038",
  1724 => x"70fd248a",
  1725 => x"3870fc2e",
  1726 => x"80cc38b6",
  1727 => x"d00470fe",
  1728 => x"2eb73870",
  1729 => x"ff2e0981",
  1730 => x"0680c538",
  1731 => x"80c0d808",
  1732 => x"5170802e",
  1733 => x"bb38ff11",
  1734 => x"80c0d80c",
  1735 => x"b6d00480",
  1736 => x"c0d808f0",
  1737 => x"057080c0",
  1738 => x"d80c5170",
  1739 => x"8025a138",
  1740 => x"800b80c0",
  1741 => x"d80cb6d0",
  1742 => x"0480c0d8",
  1743 => x"08810580",
  1744 => x"c0d80cb6",
  1745 => x"d00480c0",
  1746 => x"d8089005",
  1747 => x"80c0d80c",
  1748 => x"b2ed2d90",
  1749 => x"9d2d0284",
  1750 => x"050d0402",
  1751 => x"fc050d80",
  1752 => x"0b80c0d8",
  1753 => x"0cb2ed2d",
  1754 => x"8f9b2d80",
  1755 => x"c0dc0880",
  1756 => x"c0c80cbf",
  1757 => x"a45191bf",
  1758 => x"2d028405",
  1759 => x"0d047180",
  1760 => x"c88c0c04",
  1761 => x"00ffffff",
  1762 => x"ff00ffff",
  1763 => x"ffff00ff",
  1764 => x"ffffff00",
  1765 => x"52657365",
  1766 => x"74204e45",
  1767 => x"53000000",
  1768 => x"5363616e",
  1769 => x"6c696e65",
  1770 => x"7320284f",
  1771 => x"53442900",
  1772 => x"48713278",
  1773 => x"2066696c",
  1774 => x"74657200",
  1775 => x"466f7263",
  1776 => x"65642073",
  1777 => x"63616e64",
  1778 => x"6f75626c",
  1779 => x"65720000",
  1780 => x"48696465",
  1781 => x"206f7665",
  1782 => x"72736361",
  1783 => x"6e000000",
  1784 => x"4175746f",
  1785 => x"2d737761",
  1786 => x"702f456a",
  1787 => x"65637420",
  1788 => x"46445320",
  1789 => x"6469736b",
  1790 => x"00000000",
  1791 => x"4c6f6164",
  1792 => x"204e4553",
  1793 => x"20524f4d",
  1794 => x"20100000",
  1795 => x"4c6f6164",
  1796 => x"20506f77",
  1797 => x"65727061",
  1798 => x"6b204644",
  1799 => x"53204269",
  1800 => x"6f732010",
  1801 => x"00000000",
  1802 => x"4c6f6164",
  1803 => x"20464453",
  1804 => x"20524f4d",
  1805 => x"20100000",
  1806 => x"45786974",
  1807 => x"00000000",
  1808 => x"536d6f6f",
  1809 => x"74682070",
  1810 => x"616c6574",
  1811 => x"74650000",
  1812 => x"4e545343",
  1813 => x"20756e73",
  1814 => x"61747572",
  1815 => x"61746564",
  1816 => x"56362070",
  1817 => x"616c6574",
  1818 => x"74650000",
  1819 => x"46434555",
  1820 => x"58207061",
  1821 => x"6c657474",
  1822 => x"65000000",
  1823 => x"4e455320",
  1824 => x"636c6173",
  1825 => x"73696320",
  1826 => x"70616c65",
  1827 => x"74746500",
  1828 => x"436f6d70",
  1829 => x"6f736974",
  1830 => x"65206469",
  1831 => x"72656374",
  1832 => x"2070616c",
  1833 => x"65747465",
  1834 => x"00000000",
  1835 => x"50432d31",
  1836 => x"30207061",
  1837 => x"6c657474",
  1838 => x"65000000",
  1839 => x"50564d20",
  1840 => x"70616c65",
  1841 => x"74746500",
  1842 => x"57617665",
  1843 => x"6265616d",
  1844 => x"2070616c",
  1845 => x"65747465",
  1846 => x"00000000",
  1847 => x"5363616e",
  1848 => x"6c696e65",
  1849 => x"73206f66",
  1850 => x"66000000",
  1851 => x"5363616e",
  1852 => x"6c696e65",
  1853 => x"73203235",
  1854 => x"25000000",
  1855 => x"5363616e",
  1856 => x"6c696e65",
  1857 => x"73203530",
  1858 => x"25000000",
  1859 => x"5363616e",
  1860 => x"6c696e65",
  1861 => x"73203735",
  1862 => x"25000000",
  1863 => x"4175746f",
  1864 => x"20736964",
  1865 => x"65000000",
  1866 => x"4175746f",
  1867 => x"20736964",
  1868 => x"65202b20",
  1869 => x"31000000",
  1870 => x"4175746f",
  1871 => x"20736964",
  1872 => x"65202b20",
  1873 => x"32000000",
  1874 => x"4175746f",
  1875 => x"20736964",
  1876 => x"65202b20",
  1877 => x"33000000",
  1878 => x"524f4d20",
  1879 => x"6c6f6164",
  1880 => x"696e6720",
  1881 => x"6661696c",
  1882 => x"65640000",
  1883 => x"4f4b0000",
  1884 => x"496e6974",
  1885 => x"69616c69",
  1886 => x"7a696e67",
  1887 => x"20534420",
  1888 => x"63617264",
  1889 => x"0a000000",
  1890 => x"16200000",
  1891 => x"14200000",
  1892 => x"15200000",
  1893 => x"53442069",
  1894 => x"6e69742e",
  1895 => x"2e2e0a00",
  1896 => x"53442063",
  1897 => x"61726420",
  1898 => x"72657365",
  1899 => x"74206661",
  1900 => x"696c6564",
  1901 => x"210a0000",
  1902 => x"53444843",
  1903 => x"20657272",
  1904 => x"6f72210a",
  1905 => x"00000000",
  1906 => x"57726974",
  1907 => x"65206661",
  1908 => x"696c6564",
  1909 => x"0a000000",
  1910 => x"52656164",
  1911 => x"20666169",
  1912 => x"6c65640a",
  1913 => x"00000000",
  1914 => x"43617264",
  1915 => x"20696e69",
  1916 => x"74206661",
  1917 => x"696c6564",
  1918 => x"0a000000",
  1919 => x"46415431",
  1920 => x"36202020",
  1921 => x"00000000",
  1922 => x"46415433",
  1923 => x"32202020",
  1924 => x"00000000",
  1925 => x"4e6f2070",
  1926 => x"61727469",
  1927 => x"74696f6e",
  1928 => x"20736967",
  1929 => x"0a000000",
  1930 => x"42616420",
  1931 => x"70617274",
  1932 => x"0a000000",
  1933 => x"4261636b",
  1934 => x"00000000",
  1935 => x"00000002",
  1936 => x"00000000",
  1937 => x"00000002",
  1938 => x"00001b94",
  1939 => x"00000369",
  1940 => x"00000001",
  1941 => x"00001ba0",
  1942 => x"00000000",
  1943 => x"00000001",
  1944 => x"00001bb0",
  1945 => x"00000001",
  1946 => x"00000001",
  1947 => x"00001bbc",
  1948 => x"00000002",
  1949 => x"00000001",
  1950 => x"00001bd0",
  1951 => x"00000003",
  1952 => x"00000001",
  1953 => x"00001be0",
  1954 => x"00000004",
  1955 => x"00000003",
  1956 => x"00001f1c",
  1957 => x"00000004",
  1958 => x"00000003",
  1959 => x"00001f0c",
  1960 => x"00000004",
  1961 => x"00000003",
  1962 => x"00001eec",
  1963 => x"00000008",
  1964 => x"00000002",
  1965 => x"00001bfc",
  1966 => x"000003ae",
  1967 => x"00000002",
  1968 => x"00001c0c",
  1969 => x"000003c1",
  1970 => x"00000002",
  1971 => x"00001c28",
  1972 => x"000003d4",
  1973 => x"00000002",
  1974 => x"00001c38",
  1975 => x"000007b7",
  1976 => x"00000000",
  1977 => x"00000000",
  1978 => x"00000000",
  1979 => x"00001c40",
  1980 => x"00001c50",
  1981 => x"00001c6c",
  1982 => x"00001c7c",
  1983 => x"00001c90",
  1984 => x"00001cac",
  1985 => x"00001cbc",
  1986 => x"00001cc8",
  1987 => x"00001cdc",
  1988 => x"00001cec",
  1989 => x"00001cfc",
  1990 => x"00001d0c",
  1991 => x"00001d1c",
  1992 => x"00001d28",
  1993 => x"00001d38",
  1994 => x"00001d48",
  1995 => x"00000004",
  1996 => x"00001d58",
  1997 => x"00001f2c",
  1998 => x"00000004",
  1999 => x"00001d6c",
  2000 => x"00001e44",
  2001 => x"00000000",
  2002 => x"00000000",
  2003 => x"00000000",
  2004 => x"00000000",
  2005 => x"00000000",
  2006 => x"00000000",
  2007 => x"00000000",
  2008 => x"00000000",
  2009 => x"00000000",
  2010 => x"00000000",
  2011 => x"00000000",
  2012 => x"00000000",
  2013 => x"00000000",
  2014 => x"00000000",
  2015 => x"00000000",
  2016 => x"00000000",
  2017 => x"00000000",
  2018 => x"00000000",
  2019 => x"00000000",
  2020 => x"00000000",
  2021 => x"00000000",
  2022 => x"00000000",
  2023 => x"00000000",
  2024 => x"00000000",
  2025 => x"00000002",
  2026 => x"00002410",
  2027 => x"00001935",
  2028 => x"00000002",
  2029 => x"0000242e",
  2030 => x"00001935",
  2031 => x"00000002",
  2032 => x"0000244c",
  2033 => x"00001935",
  2034 => x"00000002",
  2035 => x"0000246a",
  2036 => x"00001935",
  2037 => x"00000002",
  2038 => x"00002488",
  2039 => x"00001935",
  2040 => x"00000002",
  2041 => x"000024a6",
  2042 => x"00001935",
  2043 => x"00000002",
  2044 => x"000024c4",
  2045 => x"00001935",
  2046 => x"00000002",
  2047 => x"000024e2",
  2048 => x"00001935",
  2049 => x"00000002",
  2050 => x"00002500",
  2051 => x"00001935",
  2052 => x"00000002",
  2053 => x"0000251e",
  2054 => x"00001935",
  2055 => x"00000002",
  2056 => x"0000253c",
  2057 => x"00001935",
  2058 => x"00000002",
  2059 => x"0000255a",
  2060 => x"00001935",
  2061 => x"00000002",
  2062 => x"00002578",
  2063 => x"00001935",
  2064 => x"00000004",
  2065 => x"00001e34",
  2066 => x"00000000",
  2067 => x"00000000",
  2068 => x"00000000",
  2069 => x"00001ae5",
  2070 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

