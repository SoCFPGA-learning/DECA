-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"0b0b0b0b",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"00000016",
     7 => x"00000000",
     8 => x"0b0b0bb8",
     9 => x"8c080b0b",
    10 => x"0bb89008",
    11 => x"0b0b0bb8",
    12 => x"94080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b0b",
    15 => x"b8940c0b",
    16 => x"0b0bb890",
    17 => x"0c0b0b0b",
    18 => x"b88c0c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b0bafdc",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"b88c7080",
    57 => x"c2bc278b",
    58 => x"38807170",
    59 => x"8405530c",
    60 => x"81e2048c",
    61 => x"51889d04",
    62 => x"02fc050d",
    63 => x"f880518f",
    64 => x"0bb89c0c",
    65 => x"9f0bb8a0",
    66 => x"0ca07170",
    67 => x"81055334",
    68 => x"b8a008ff",
    69 => x"05b8a00c",
    70 => x"b8a00880",
    71 => x"25eb38b8",
    72 => x"9c08ff05",
    73 => x"b89c0cb8",
    74 => x"9c088025",
    75 => x"d738800b",
    76 => x"b8a00c80",
    77 => x"0bb89c0c",
    78 => x"0284050d",
    79 => x"0402f005",
    80 => x"0df88053",
    81 => x"f8a05483",
    82 => x"bf527370",
    83 => x"81055533",
    84 => x"51707370",
    85 => x"81055534",
    86 => x"ff125271",
    87 => x"8025eb38",
    88 => x"fbc0539f",
    89 => x"52a07370",
    90 => x"81055534",
    91 => x"ff125271",
    92 => x"8025f238",
    93 => x"0290050d",
    94 => x"0402f405",
    95 => x"0d74538e",
    96 => x"0bb89c08",
    97 => x"258f3882",
    98 => x"bd2db89c",
    99 => x"08ff05b8",
   100 => x"9c0c82ff",
   101 => x"04b89c08",
   102 => x"b8a00853",
   103 => x"51728a2e",
   104 => x"098106b7",
   105 => x"38715171",
   106 => x"9f24a038",
   107 => x"b89c08a0",
   108 => x"2911f880",
   109 => x"115151a0",
   110 => x"7134b8a0",
   111 => x"088105b8",
   112 => x"a00cb8a0",
   113 => x"08519f71",
   114 => x"25e23880",
   115 => x"0bb8a00c",
   116 => x"b89c0881",
   117 => x"05b89c0c",
   118 => x"83ef0470",
   119 => x"a02912f8",
   120 => x"80115151",
   121 => x"727134b8",
   122 => x"a0088105",
   123 => x"b8a00cb8",
   124 => x"a008a02e",
   125 => x"0981068e",
   126 => x"38800bb8",
   127 => x"a00cb89c",
   128 => x"088105b8",
   129 => x"9c0c028c",
   130 => x"050d0402",
   131 => x"e8050d77",
   132 => x"79565688",
   133 => x"0bfc1677",
   134 => x"712c8f06",
   135 => x"54525480",
   136 => x"53727225",
   137 => x"95387153",
   138 => x"fbe01451",
   139 => x"87713481",
   140 => x"14ff1454",
   141 => x"5472f138",
   142 => x"7153f915",
   143 => x"76712c87",
   144 => x"06535171",
   145 => x"802e8b38",
   146 => x"fbe01451",
   147 => x"71713481",
   148 => x"1454728e",
   149 => x"2495388f",
   150 => x"733153fb",
   151 => x"e01451a0",
   152 => x"71348114",
   153 => x"ff145454",
   154 => x"72f13802",
   155 => x"98050d04",
   156 => x"02ec050d",
   157 => x"800bb8a4",
   158 => x"0cf68c08",
   159 => x"f6900871",
   160 => x"882c5654",
   161 => x"81ff0652",
   162 => x"73722588",
   163 => x"38715482",
   164 => x"0bb8a40c",
   165 => x"72882c73",
   166 => x"81ff0654",
   167 => x"55747325",
   168 => x"8b3872b8",
   169 => x"a4088407",
   170 => x"b8a40c55",
   171 => x"73842b86",
   172 => x"a0712583",
   173 => x"7131700b",
   174 => x"0b0bb490",
   175 => x"0c81712b",
   176 => x"ff05f688",
   177 => x"0cfdfc13",
   178 => x"ff122c78",
   179 => x"8829ff94",
   180 => x"0570812c",
   181 => x"b8a40852",
   182 => x"58525551",
   183 => x"52547680",
   184 => x"2e853870",
   185 => x"81075170",
   186 => x"f6940c71",
   187 => x"098105f6",
   188 => x"800c7209",
   189 => x"8105f684",
   190 => x"0c029405",
   191 => x"0d0402f4",
   192 => x"050d7453",
   193 => x"72708105",
   194 => x"5480f52d",
   195 => x"5271802e",
   196 => x"89387151",
   197 => x"82f92d86",
   198 => x"8404810b",
   199 => x"b88c0c02",
   200 => x"8c050d04",
   201 => x"02fc050d",
   202 => x"81808051",
   203 => x"c0115170",
   204 => x"fb380284",
   205 => x"050d0402",
   206 => x"fc050d84",
   207 => x"bf5186a4",
   208 => x"2dff1151",
   209 => x"708025f6",
   210 => x"38028405",
   211 => x"0d0402fc",
   212 => x"050dec51",
   213 => x"83710c86",
   214 => x"a42d8271",
   215 => x"0c028405",
   216 => x"0d04880b",
   217 => x"ec0c86b7",
   218 => x"2d0402dc",
   219 => x"050d8059",
   220 => x"86e22d90",
   221 => x"0bec0c7a",
   222 => x"52b8a851",
   223 => x"a7982db8",
   224 => x"8c08792e",
   225 => x"80ee38b8",
   226 => x"ac0870f8",
   227 => x"0c79ff12",
   228 => x"56595573",
   229 => x"792e8b38",
   230 => x"81187481",
   231 => x"2a555873",
   232 => x"f738f718",
   233 => x"58815980",
   234 => x"752580c8",
   235 => x"38775273",
   236 => x"51848b2d",
   237 => x"b8f452b8",
   238 => x"a851a9ce",
   239 => x"2db88c08",
   240 => x"802e9a38",
   241 => x"b8f45783",
   242 => x"fc567670",
   243 => x"84055808",
   244 => x"e80cfc16",
   245 => x"56758025",
   246 => x"f13887e4",
   247 => x"04b88c08",
   248 => x"59848055",
   249 => x"b8a851a9",
   250 => x"a12dfc80",
   251 => x"15811555",
   252 => x"5587a704",
   253 => x"805186ce",
   254 => x"2d840bec",
   255 => x"0c78802e",
   256 => x"8d38b494",
   257 => x"5190a62d",
   258 => x"8ea92d88",
   259 => x"9404b5dc",
   260 => x"5190a62d",
   261 => x"78b88c0c",
   262 => x"02a4050d",
   263 => x"0402ec05",
   264 => x"0d840bec",
   265 => x"0c8df72d",
   266 => x"8ac62d81",
   267 => x"f82d8352",
   268 => x"8ddc2d81",
   269 => x"5184f02d",
   270 => x"ff125271",
   271 => x"8025f138",
   272 => x"840bec0c",
   273 => x"b2c45185",
   274 => x"fe2d9eb5",
   275 => x"2db88c08",
   276 => x"802e81dd",
   277 => x"3886ea51",
   278 => x"afd52db4",
   279 => x"945190a6",
   280 => x"2d8e962d",
   281 => x"8ad22d90",
   282 => x"b62db88c",
   283 => x"08b4c00b",
   284 => x"80f52db6",
   285 => x"c8087081",
   286 => x"06555654",
   287 => x"5571802e",
   288 => x"85387284",
   289 => x"07537381",
   290 => x"2a708106",
   291 => x"51527180",
   292 => x"2e853872",
   293 => x"88075373",
   294 => x"822a7081",
   295 => x"06515271",
   296 => x"802e8538",
   297 => x"72900753",
   298 => x"73832a70",
   299 => x"81065152",
   300 => x"71802e85",
   301 => x"3872a007",
   302 => x"53b4e40b",
   303 => x"80f52d52",
   304 => x"71812e09",
   305 => x"81068938",
   306 => x"7280c007",
   307 => x"5389ed04",
   308 => x"71822e09",
   309 => x"81068938",
   310 => x"72818007",
   311 => x"5389ed04",
   312 => x"71832e09",
   313 => x"81068638",
   314 => x"7281c007",
   315 => x"53b4f00b",
   316 => x"80f52d52",
   317 => x"71812e09",
   318 => x"81068938",
   319 => x"72828007",
   320 => x"538aa104",
   321 => x"71822e09",
   322 => x"81068938",
   323 => x"72848007",
   324 => x"538aa104",
   325 => x"71832e09",
   326 => x"81068638",
   327 => x"72868007",
   328 => x"5372fc0c",
   329 => x"86527483",
   330 => x"38845271",
   331 => x"ec0c88e4",
   332 => x"04800bb8",
   333 => x"8c0c0294",
   334 => x"050d0471",
   335 => x"980c04ff",
   336 => x"b008b88c",
   337 => x"0c04810b",
   338 => x"ffb00c04",
   339 => x"800bffb0",
   340 => x"0c0402f4",
   341 => x"050d8bd4",
   342 => x"04b88c08",
   343 => x"81f02e09",
   344 => x"81068938",
   345 => x"810bb6c0",
   346 => x"0c8bd404",
   347 => x"b88c0881",
   348 => x"e02e0981",
   349 => x"06893881",
   350 => x"0bb6c40c",
   351 => x"8bd404b8",
   352 => x"8c0852b6",
   353 => x"c408802e",
   354 => x"8838b88c",
   355 => x"08818005",
   356 => x"5271842c",
   357 => x"728f0653",
   358 => x"53b6c008",
   359 => x"802e9938",
   360 => x"728429b6",
   361 => x"80057213",
   362 => x"81712b70",
   363 => x"09730806",
   364 => x"730c5153",
   365 => x"538bca04",
   366 => x"728429b6",
   367 => x"80057213",
   368 => x"83712b72",
   369 => x"0807720c",
   370 => x"5353800b",
   371 => x"b6c40c80",
   372 => x"0bb6c00c",
   373 => x"b8b4518c",
   374 => x"d52db88c",
   375 => x"08ff24fe",
   376 => x"f838800b",
   377 => x"b88c0c02",
   378 => x"8c050d04",
   379 => x"02f8050d",
   380 => x"b680528f",
   381 => x"51807270",
   382 => x"8405540c",
   383 => x"ff115170",
   384 => x"8025f238",
   385 => x"0288050d",
   386 => x"0402f005",
   387 => x"0d75518a",
   388 => x"cc2d7082",
   389 => x"2cfc06b6",
   390 => x"80117210",
   391 => x"9e067108",
   392 => x"70722a70",
   393 => x"83068274",
   394 => x"2b700974",
   395 => x"06760c54",
   396 => x"51565753",
   397 => x"51538ac6",
   398 => x"2d71b88c",
   399 => x"0c029005",
   400 => x"0d0402fc",
   401 => x"050d7251",
   402 => x"80710c80",
   403 => x"0b84120c",
   404 => x"0284050d",
   405 => x"0402f005",
   406 => x"0d757008",
   407 => x"84120853",
   408 => x"5353ff54",
   409 => x"71712ea8",
   410 => x"388acc2d",
   411 => x"84130870",
   412 => x"84291488",
   413 => x"11700870",
   414 => x"81ff0684",
   415 => x"18088111",
   416 => x"8706841a",
   417 => x"0c535155",
   418 => x"5151518a",
   419 => x"c62d7154",
   420 => x"73b88c0c",
   421 => x"0290050d",
   422 => x"0402f805",
   423 => x"0d8acc2d",
   424 => x"e008708b",
   425 => x"2a708106",
   426 => x"51525270",
   427 => x"802e9d38",
   428 => x"b8b40870",
   429 => x"8429b8bc",
   430 => x"057381ff",
   431 => x"06710c51",
   432 => x"51b8b408",
   433 => x"81118706",
   434 => x"b8b40c51",
   435 => x"800bb8dc",
   436 => x"0c8abf2d",
   437 => x"8ac62d02",
   438 => x"88050d04",
   439 => x"02fc050d",
   440 => x"8acc2d81",
   441 => x"0bb8dc0c",
   442 => x"8ac62db8",
   443 => x"dc085170",
   444 => x"fa380284",
   445 => x"050d0402",
   446 => x"fc050db8",
   447 => x"b4518cc2",
   448 => x"2d8bec2d",
   449 => x"8d99518a",
   450 => x"bb2d0284",
   451 => x"050d04b8",
   452 => x"e008b88c",
   453 => x"0c0402fc",
   454 => x"050d810b",
   455 => x"b6cc0c81",
   456 => x"5184f02d",
   457 => x"0284050d",
   458 => x"0402fc05",
   459 => x"0d8eb304",
   460 => x"8ad22d80",
   461 => x"f6518c89",
   462 => x"2db88c08",
   463 => x"f33880da",
   464 => x"518c892d",
   465 => x"b88c08e8",
   466 => x"38b88c08",
   467 => x"b6cc0cb8",
   468 => x"8c085184",
   469 => x"f02d0284",
   470 => x"050d0402",
   471 => x"ec050d76",
   472 => x"54805287",
   473 => x"0b881580",
   474 => x"f52d5653",
   475 => x"74722483",
   476 => x"38a05372",
   477 => x"5182f92d",
   478 => x"81128b15",
   479 => x"80f52d54",
   480 => x"52727225",
   481 => x"de380294",
   482 => x"050d0402",
   483 => x"f0050db8",
   484 => x"e0085481",
   485 => x"f82d800b",
   486 => x"b8e40c73",
   487 => x"08802e81",
   488 => x"8038820b",
   489 => x"b8a00cb8",
   490 => x"e4088f06",
   491 => x"b89c0c73",
   492 => x"08527183",
   493 => x"2e963871",
   494 => x"83268938",
   495 => x"71812eaf",
   496 => x"38908c04",
   497 => x"71852e9f",
   498 => x"38908c04",
   499 => x"881480f5",
   500 => x"2d841508",
   501 => x"b2dc5354",
   502 => x"5285fe2d",
   503 => x"71842913",
   504 => x"70085252",
   505 => x"90900473",
   506 => x"518edb2d",
   507 => x"908c04b6",
   508 => x"c8088815",
   509 => x"082c7081",
   510 => x"06515271",
   511 => x"802e8738",
   512 => x"b2e05190",
   513 => x"8904b2e4",
   514 => x"5185fe2d",
   515 => x"84140851",
   516 => x"85fe2db8",
   517 => x"e4088105",
   518 => x"b8e40c8c",
   519 => x"14548f9b",
   520 => x"04029005",
   521 => x"0d0471b8",
   522 => x"e00c8f8b",
   523 => x"2db8e408",
   524 => x"ff05b8e8",
   525 => x"0c0402e8",
   526 => x"050db8e0",
   527 => x"08b8ec08",
   528 => x"575580f6",
   529 => x"518c892d",
   530 => x"b88c0881",
   531 => x"2a708106",
   532 => x"51527180",
   533 => x"2ea13890",
   534 => x"dd048ad2",
   535 => x"2d80f651",
   536 => x"8c892db8",
   537 => x"8c08f338",
   538 => x"b6cc0881",
   539 => x"3270b6cc",
   540 => x"0c705252",
   541 => x"84f02db6",
   542 => x"cc089038",
   543 => x"81fd518c",
   544 => x"892d81fa",
   545 => x"518c892d",
   546 => x"96bc0481",
   547 => x"f5518c89",
   548 => x"2db88c08",
   549 => x"812a7081",
   550 => x"06515271",
   551 => x"802eaf38",
   552 => x"b8e80852",
   553 => x"71802e89",
   554 => x"38ff12b8",
   555 => x"e80c91ce",
   556 => x"04b8e408",
   557 => x"10b8e408",
   558 => x"05708429",
   559 => x"16515288",
   560 => x"1208802e",
   561 => x"8938ff51",
   562 => x"88120852",
   563 => x"712d81f2",
   564 => x"518c892d",
   565 => x"b88c0881",
   566 => x"2a708106",
   567 => x"51527180",
   568 => x"2eb138b8",
   569 => x"e408ff11",
   570 => x"b8e80856",
   571 => x"53537372",
   572 => x"25893881",
   573 => x"14b8e80c",
   574 => x"92930472",
   575 => x"10137084",
   576 => x"29165152",
   577 => x"88120880",
   578 => x"2e8938fe",
   579 => x"51881208",
   580 => x"52712d81",
   581 => x"fd518c89",
   582 => x"2db88c08",
   583 => x"812a7081",
   584 => x"06515271",
   585 => x"802ead38",
   586 => x"b8e80880",
   587 => x"2e893880",
   588 => x"0bb8e80c",
   589 => x"92d404b8",
   590 => x"e40810b8",
   591 => x"e4080570",
   592 => x"84291651",
   593 => x"52881208",
   594 => x"802e8938",
   595 => x"fd518812",
   596 => x"0852712d",
   597 => x"81fa518c",
   598 => x"892db88c",
   599 => x"08812a70",
   600 => x"81065152",
   601 => x"71802eae",
   602 => x"38b8e408",
   603 => x"ff115452",
   604 => x"b8e80873",
   605 => x"25883872",
   606 => x"b8e80c93",
   607 => x"96047110",
   608 => x"12708429",
   609 => x"16515288",
   610 => x"1208802e",
   611 => x"8938fc51",
   612 => x"88120852",
   613 => x"712db8e8",
   614 => x"08705354",
   615 => x"73802e8a",
   616 => x"388c15ff",
   617 => x"15555593",
   618 => x"9c04820b",
   619 => x"b8a00c71",
   620 => x"8f06b89c",
   621 => x"0c81eb51",
   622 => x"8c892db8",
   623 => x"8c08812a",
   624 => x"70810651",
   625 => x"5271802e",
   626 => x"ad387408",
   627 => x"852e0981",
   628 => x"06a43888",
   629 => x"1580f52d",
   630 => x"ff055271",
   631 => x"881681b7",
   632 => x"2d71982b",
   633 => x"52718025",
   634 => x"8838800b",
   635 => x"881681b7",
   636 => x"2d74518e",
   637 => x"db2d81f4",
   638 => x"518c892d",
   639 => x"b88c0881",
   640 => x"2a708106",
   641 => x"51527180",
   642 => x"2eb33874",
   643 => x"08852e09",
   644 => x"8106aa38",
   645 => x"881580f5",
   646 => x"2d810552",
   647 => x"71881681",
   648 => x"b72d7181",
   649 => x"ff068b16",
   650 => x"80f52d54",
   651 => x"52727227",
   652 => x"87387288",
   653 => x"1681b72d",
   654 => x"74518edb",
   655 => x"2d80da51",
   656 => x"8c892db8",
   657 => x"8c08812a",
   658 => x"70810651",
   659 => x"5271802e",
   660 => x"81a638b8",
   661 => x"e008b8e8",
   662 => x"08555373",
   663 => x"802e8a38",
   664 => x"8c13ff15",
   665 => x"555394db",
   666 => x"04720852",
   667 => x"71822ea6",
   668 => x"38718226",
   669 => x"89387181",
   670 => x"2ea93895",
   671 => x"f8047183",
   672 => x"2eb13871",
   673 => x"842e0981",
   674 => x"0680ed38",
   675 => x"88130851",
   676 => x"90a62d95",
   677 => x"f804b8e8",
   678 => x"08518813",
   679 => x"0852712d",
   680 => x"95f80481",
   681 => x"0b881408",
   682 => x"2bb6c808",
   683 => x"32b6c80c",
   684 => x"95ce0488",
   685 => x"1380f52d",
   686 => x"81058b14",
   687 => x"80f52d53",
   688 => x"54717424",
   689 => x"83388054",
   690 => x"73881481",
   691 => x"b72d8f8b",
   692 => x"2d95f804",
   693 => x"7508802e",
   694 => x"a2387508",
   695 => x"518c892d",
   696 => x"b88c0881",
   697 => x"06527180",
   698 => x"2e8b38b8",
   699 => x"e8085184",
   700 => x"16085271",
   701 => x"2d881656",
   702 => x"75da3880",
   703 => x"54800bb8",
   704 => x"a00c738f",
   705 => x"06b89c0c",
   706 => x"a05273b8",
   707 => x"e8082e09",
   708 => x"81069838",
   709 => x"b8e408ff",
   710 => x"05743270",
   711 => x"09810570",
   712 => x"72079f2a",
   713 => x"91713151",
   714 => x"51535371",
   715 => x"5182f92d",
   716 => x"8114548e",
   717 => x"7425c638",
   718 => x"b6cc0852",
   719 => x"71b88c0c",
   720 => x"0298050d",
   721 => x"0402f405",
   722 => x"0dd45281",
   723 => x"ff720c71",
   724 => x"085381ff",
   725 => x"720c7288",
   726 => x"2b83fe80",
   727 => x"06720870",
   728 => x"81ff0651",
   729 => x"525381ff",
   730 => x"720c7271",
   731 => x"07882b72",
   732 => x"087081ff",
   733 => x"06515253",
   734 => x"81ff720c",
   735 => x"72710788",
   736 => x"2b720870",
   737 => x"81ff0672",
   738 => x"07b88c0c",
   739 => x"5253028c",
   740 => x"050d0402",
   741 => x"f4050d74",
   742 => x"767181ff",
   743 => x"06d40c53",
   744 => x"53b8f008",
   745 => x"85387189",
   746 => x"2b527198",
   747 => x"2ad40c71",
   748 => x"902a7081",
   749 => x"ff06d40c",
   750 => x"5171882a",
   751 => x"7081ff06",
   752 => x"d40c5171",
   753 => x"81ff06d4",
   754 => x"0c72902a",
   755 => x"7081ff06",
   756 => x"d40c51d4",
   757 => x"087081ff",
   758 => x"06515182",
   759 => x"b8bf5270",
   760 => x"81ff2e09",
   761 => x"81069438",
   762 => x"81ff0bd4",
   763 => x"0cd40870",
   764 => x"81ff06ff",
   765 => x"14545151",
   766 => x"71e53870",
   767 => x"b88c0c02",
   768 => x"8c050d04",
   769 => x"02fc050d",
   770 => x"81c75181",
   771 => x"ff0bd40c",
   772 => x"ff115170",
   773 => x"8025f438",
   774 => x"0284050d",
   775 => x"0402f405",
   776 => x"0d81ff0b",
   777 => x"d40c9353",
   778 => x"805287fc",
   779 => x"80c15197",
   780 => x"932db88c",
   781 => x"088b3881",
   782 => x"ff0bd40c",
   783 => x"815398ca",
   784 => x"0498842d",
   785 => x"ff135372",
   786 => x"df3872b8",
   787 => x"8c0c028c",
   788 => x"050d0402",
   789 => x"ec050d81",
   790 => x"0bb8f00c",
   791 => x"8454d008",
   792 => x"708f2a70",
   793 => x"81065151",
   794 => x"5372f338",
   795 => x"72d00c98",
   796 => x"842db2e8",
   797 => x"5185fe2d",
   798 => x"d008708f",
   799 => x"2a708106",
   800 => x"51515372",
   801 => x"f338810b",
   802 => x"d00cb153",
   803 => x"805284d4",
   804 => x"80c05197",
   805 => x"932db88c",
   806 => x"08812e93",
   807 => x"3872822e",
   808 => x"bd38ff13",
   809 => x"5372e538",
   810 => x"ff145473",
   811 => x"ffb03898",
   812 => x"842d83aa",
   813 => x"52849c80",
   814 => x"c8519793",
   815 => x"2db88c08",
   816 => x"812e0981",
   817 => x"06923896",
   818 => x"c52db88c",
   819 => x"0883ffff",
   820 => x"06537283",
   821 => x"aa2e9d38",
   822 => x"989d2d99",
   823 => x"ef04b2f4",
   824 => x"5185fe2d",
   825 => x"80539bbd",
   826 => x"04b38c51",
   827 => x"85fe2d80",
   828 => x"549b8f04",
   829 => x"81ff0bd4",
   830 => x"0cb15498",
   831 => x"842d8fcf",
   832 => x"53805287",
   833 => x"fc80f751",
   834 => x"97932db8",
   835 => x"8c0855b8",
   836 => x"8c08812e",
   837 => x"0981069b",
   838 => x"3881ff0b",
   839 => x"d40c820a",
   840 => x"52849c80",
   841 => x"e9519793",
   842 => x"2db88c08",
   843 => x"802e8d38",
   844 => x"98842dff",
   845 => x"135372c9",
   846 => x"389b8204",
   847 => x"81ff0bd4",
   848 => x"0cb88c08",
   849 => x"5287fc80",
   850 => x"fa519793",
   851 => x"2db88c08",
   852 => x"b13881ff",
   853 => x"0bd40cd4",
   854 => x"085381ff",
   855 => x"0bd40c81",
   856 => x"ff0bd40c",
   857 => x"81ff0bd4",
   858 => x"0c81ff0b",
   859 => x"d40c7286",
   860 => x"2a708106",
   861 => x"76565153",
   862 => x"729538b8",
   863 => x"8c08549b",
   864 => x"8f047382",
   865 => x"2efee238",
   866 => x"ff145473",
   867 => x"feed3873",
   868 => x"b8f00c73",
   869 => x"8b388152",
   870 => x"87fc80d0",
   871 => x"5197932d",
   872 => x"81ff0bd4",
   873 => x"0cd00870",
   874 => x"8f2a7081",
   875 => x"06515153",
   876 => x"72f33872",
   877 => x"d00c81ff",
   878 => x"0bd40c81",
   879 => x"5372b88c",
   880 => x"0c029405",
   881 => x"0d0402e8",
   882 => x"050d7855",
   883 => x"805681ff",
   884 => x"0bd40cd0",
   885 => x"08708f2a",
   886 => x"70810651",
   887 => x"515372f3",
   888 => x"3882810b",
   889 => x"d00c81ff",
   890 => x"0bd40c77",
   891 => x"5287fc80",
   892 => x"d1519793",
   893 => x"2d80dbc6",
   894 => x"df54b88c",
   895 => x"08802e8a",
   896 => x"38b3ac51",
   897 => x"85fe2d9c",
   898 => x"dd0481ff",
   899 => x"0bd40cd4",
   900 => x"087081ff",
   901 => x"06515372",
   902 => x"81fe2e09",
   903 => x"81069d38",
   904 => x"80ff5396",
   905 => x"c52db88c",
   906 => x"08757084",
   907 => x"05570cff",
   908 => x"13537280",
   909 => x"25ed3881",
   910 => x"569cc204",
   911 => x"ff145473",
   912 => x"c93881ff",
   913 => x"0bd40c81",
   914 => x"ff0bd40c",
   915 => x"d008708f",
   916 => x"2a708106",
   917 => x"51515372",
   918 => x"f33872d0",
   919 => x"0c75b88c",
   920 => x"0c029805",
   921 => x"0d0402e8",
   922 => x"050d7779",
   923 => x"7b585555",
   924 => x"80537276",
   925 => x"25a33874",
   926 => x"70810556",
   927 => x"80f52d74",
   928 => x"70810556",
   929 => x"80f52d52",
   930 => x"5271712e",
   931 => x"86388151",
   932 => x"9d9b0481",
   933 => x"13539cf2",
   934 => x"04805170",
   935 => x"b88c0c02",
   936 => x"98050d04",
   937 => x"02ec050d",
   938 => x"76557480",
   939 => x"2ebb389a",
   940 => x"1580e02d",
   941 => x"51aaa42d",
   942 => x"b88c08b8",
   943 => x"8c08bfa4",
   944 => x"0cb88c08",
   945 => x"5454bf80",
   946 => x"08802e99",
   947 => x"38941580",
   948 => x"e02d51aa",
   949 => x"a42db88c",
   950 => x"08902b83",
   951 => x"fff00a06",
   952 => x"70750751",
   953 => x"5372bfa4",
   954 => x"0cbfa408",
   955 => x"5372802e",
   956 => x"9938bef8",
   957 => x"08fe1471",
   958 => x"29bf8c08",
   959 => x"05bfa80c",
   960 => x"70842bbf",
   961 => x"840c549e",
   962 => x"b004bf90",
   963 => x"08bfa40c",
   964 => x"bf9408bf",
   965 => x"a80cbf80",
   966 => x"08802e8a",
   967 => x"38bef808",
   968 => x"842b539e",
   969 => x"ac04bf98",
   970 => x"08842b53",
   971 => x"72bf840c",
   972 => x"0294050d",
   973 => x"0402d805",
   974 => x"0d800bbf",
   975 => x"800c8454",
   976 => x"98d32db8",
   977 => x"8c08802e",
   978 => x"9538b8f4",
   979 => x"5280519b",
   980 => x"c62db88c",
   981 => x"08802e86",
   982 => x"38fe549e",
   983 => x"e604ff14",
   984 => x"54738024",
   985 => x"db38738c",
   986 => x"38b3bc51",
   987 => x"85fe2d73",
   988 => x"55a3ef04",
   989 => x"8056810b",
   990 => x"bfac0c88",
   991 => x"53b3d052",
   992 => x"b9aa519c",
   993 => x"e62db88c",
   994 => x"08762e09",
   995 => x"81068738",
   996 => x"b88c08bf",
   997 => x"ac0c8853",
   998 => x"b3dc52b9",
   999 => x"c6519ce6",
  1000 => x"2db88c08",
  1001 => x"8738b88c",
  1002 => x"08bfac0c",
  1003 => x"bfac0880",
  1004 => x"2e80f638",
  1005 => x"bcba0b80",
  1006 => x"f52dbcbb",
  1007 => x"0b80f52d",
  1008 => x"71982b71",
  1009 => x"902b07bc",
  1010 => x"bc0b80f5",
  1011 => x"2d70882b",
  1012 => x"7207bcbd",
  1013 => x"0b80f52d",
  1014 => x"7107bcf2",
  1015 => x"0b80f52d",
  1016 => x"bcf30b80",
  1017 => x"f52d7188",
  1018 => x"2b07535f",
  1019 => x"54525a56",
  1020 => x"57557381",
  1021 => x"abaa2e09",
  1022 => x"81068d38",
  1023 => x"7551a9f4",
  1024 => x"2db88c08",
  1025 => x"56a09504",
  1026 => x"7382d4d5",
  1027 => x"2e8738b3",
  1028 => x"e851a0d6",
  1029 => x"04b8f452",
  1030 => x"75519bc6",
  1031 => x"2db88c08",
  1032 => x"55b88c08",
  1033 => x"802e83c7",
  1034 => x"388853b3",
  1035 => x"dc52b9c6",
  1036 => x"519ce62d",
  1037 => x"b88c0889",
  1038 => x"38810bbf",
  1039 => x"800ca0dc",
  1040 => x"048853b3",
  1041 => x"d052b9aa",
  1042 => x"519ce62d",
  1043 => x"b88c0880",
  1044 => x"2e8a38b3",
  1045 => x"fc5185fe",
  1046 => x"2da1b604",
  1047 => x"bcf20b80",
  1048 => x"f52d5473",
  1049 => x"80d52e09",
  1050 => x"810680ca",
  1051 => x"38bcf30b",
  1052 => x"80f52d54",
  1053 => x"7381aa2e",
  1054 => x"098106ba",
  1055 => x"38800bb8",
  1056 => x"f40b80f5",
  1057 => x"2d565474",
  1058 => x"81e92e83",
  1059 => x"38815474",
  1060 => x"81eb2e8c",
  1061 => x"38805573",
  1062 => x"752e0981",
  1063 => x"0682d038",
  1064 => x"b8ff0b80",
  1065 => x"f52d5574",
  1066 => x"8d38b980",
  1067 => x"0b80f52d",
  1068 => x"5473822e",
  1069 => x"86388055",
  1070 => x"a3ef04b9",
  1071 => x"810b80f5",
  1072 => x"2d70bef8",
  1073 => x"0cff05be",
  1074 => x"fc0cb982",
  1075 => x"0b80f52d",
  1076 => x"b9830b80",
  1077 => x"f52d5876",
  1078 => x"05778280",
  1079 => x"290570bf",
  1080 => x"880cb984",
  1081 => x"0b80f52d",
  1082 => x"70bf9c0c",
  1083 => x"bf800859",
  1084 => x"57587680",
  1085 => x"2e81a338",
  1086 => x"8853b3dc",
  1087 => x"52b9c651",
  1088 => x"9ce62db8",
  1089 => x"8c0881e7",
  1090 => x"38bef808",
  1091 => x"70842bbf",
  1092 => x"840c70bf",
  1093 => x"980cb999",
  1094 => x"0b80f52d",
  1095 => x"b9980b80",
  1096 => x"f52d7182",
  1097 => x"802905b9",
  1098 => x"9a0b80f5",
  1099 => x"2d708480",
  1100 => x"802912b9",
  1101 => x"9b0b80f5",
  1102 => x"2d708180",
  1103 => x"0a291270",
  1104 => x"bfa00cbf",
  1105 => x"9c087129",
  1106 => x"bf880805",
  1107 => x"70bf8c0c",
  1108 => x"b9a10b80",
  1109 => x"f52db9a0",
  1110 => x"0b80f52d",
  1111 => x"71828029",
  1112 => x"05b9a20b",
  1113 => x"80f52d70",
  1114 => x"84808029",
  1115 => x"12b9a30b",
  1116 => x"80f52d70",
  1117 => x"982b81f0",
  1118 => x"0a067205",
  1119 => x"70bf900c",
  1120 => x"fe117e29",
  1121 => x"7705bf94",
  1122 => x"0c525952",
  1123 => x"43545e51",
  1124 => x"5259525d",
  1125 => x"575957a3",
  1126 => x"e804b986",
  1127 => x"0b80f52d",
  1128 => x"b9850b80",
  1129 => x"f52d7182",
  1130 => x"80290570",
  1131 => x"bf840c70",
  1132 => x"a02983ff",
  1133 => x"0570892a",
  1134 => x"70bf980c",
  1135 => x"b98b0b80",
  1136 => x"f52db98a",
  1137 => x"0b80f52d",
  1138 => x"71828029",
  1139 => x"0570bfa0",
  1140 => x"0c7b7129",
  1141 => x"1e70bf94",
  1142 => x"0c7dbf90",
  1143 => x"0c7305bf",
  1144 => x"8c0c555e",
  1145 => x"51515555",
  1146 => x"80519da4",
  1147 => x"2d815574",
  1148 => x"b88c0c02",
  1149 => x"a8050d04",
  1150 => x"02ec050d",
  1151 => x"7670872c",
  1152 => x"7180ff06",
  1153 => x"555654bf",
  1154 => x"80088a38",
  1155 => x"73882c74",
  1156 => x"81ff0654",
  1157 => x"55b8f452",
  1158 => x"bf880815",
  1159 => x"519bc62d",
  1160 => x"b88c0854",
  1161 => x"b88c0880",
  1162 => x"2eb338bf",
  1163 => x"8008802e",
  1164 => x"98387284",
  1165 => x"29b8f405",
  1166 => x"70085253",
  1167 => x"a9f42db8",
  1168 => x"8c08f00a",
  1169 => x"0653a4db",
  1170 => x"047210b8",
  1171 => x"f4057080",
  1172 => x"e02d5253",
  1173 => x"aaa42db8",
  1174 => x"8c085372",
  1175 => x"5473b88c",
  1176 => x"0c029405",
  1177 => x"0d0402e0",
  1178 => x"050d7970",
  1179 => x"842cbfa8",
  1180 => x"0805718f",
  1181 => x"06525553",
  1182 => x"728938b8",
  1183 => x"f4527351",
  1184 => x"9bc62d72",
  1185 => x"a029b8f4",
  1186 => x"05548074",
  1187 => x"80f52d56",
  1188 => x"5374732e",
  1189 => x"83388153",
  1190 => x"7481e52e",
  1191 => x"81ef3881",
  1192 => x"70740654",
  1193 => x"5872802e",
  1194 => x"81e3388b",
  1195 => x"1480f52d",
  1196 => x"70832a79",
  1197 => x"06585676",
  1198 => x"9838b6d0",
  1199 => x"08537288",
  1200 => x"3872bcf4",
  1201 => x"0b81b72d",
  1202 => x"76b6d00c",
  1203 => x"7353a78f",
  1204 => x"04758f2e",
  1205 => x"09810681",
  1206 => x"b438749f",
  1207 => x"068d29bc",
  1208 => x"e7115153",
  1209 => x"811480f5",
  1210 => x"2d737081",
  1211 => x"055581b7",
  1212 => x"2d831480",
  1213 => x"f52d7370",
  1214 => x"81055581",
  1215 => x"b72d8514",
  1216 => x"80f52d73",
  1217 => x"70810555",
  1218 => x"81b72d87",
  1219 => x"1480f52d",
  1220 => x"73708105",
  1221 => x"5581b72d",
  1222 => x"891480f5",
  1223 => x"2d737081",
  1224 => x"055581b7",
  1225 => x"2d8e1480",
  1226 => x"f52d7370",
  1227 => x"81055581",
  1228 => x"b72d9014",
  1229 => x"80f52d73",
  1230 => x"70810555",
  1231 => x"81b72d92",
  1232 => x"1480f52d",
  1233 => x"73708105",
  1234 => x"5581b72d",
  1235 => x"941480f5",
  1236 => x"2d737081",
  1237 => x"055581b7",
  1238 => x"2d961480",
  1239 => x"f52d7370",
  1240 => x"81055581",
  1241 => x"b72d9814",
  1242 => x"80f52d73",
  1243 => x"70810555",
  1244 => x"81b72d9c",
  1245 => x"1480f52d",
  1246 => x"73708105",
  1247 => x"5581b72d",
  1248 => x"9e1480f5",
  1249 => x"2d7381b7",
  1250 => x"2d77b6d0",
  1251 => x"0c805372",
  1252 => x"b88c0c02",
  1253 => x"a0050d04",
  1254 => x"02cc050d",
  1255 => x"7e605e5a",
  1256 => x"800bbfa4",
  1257 => x"08bfa808",
  1258 => x"595c5680",
  1259 => x"58bf8408",
  1260 => x"782e81ae",
  1261 => x"38778f06",
  1262 => x"a0175754",
  1263 => x"738f38b8",
  1264 => x"f4527651",
  1265 => x"8117579b",
  1266 => x"c62db8f4",
  1267 => x"56807680",
  1268 => x"f52d5654",
  1269 => x"74742e83",
  1270 => x"38815474",
  1271 => x"81e52e80",
  1272 => x"f6388170",
  1273 => x"7506555c",
  1274 => x"73802e80",
  1275 => x"ea388b16",
  1276 => x"80f52d98",
  1277 => x"06597880",
  1278 => x"de388b53",
  1279 => x"7c527551",
  1280 => x"9ce62db8",
  1281 => x"8c0880cf",
  1282 => x"389c1608",
  1283 => x"51a9f42d",
  1284 => x"b88c0884",
  1285 => x"1b0c9a16",
  1286 => x"80e02d51",
  1287 => x"aaa42db8",
  1288 => x"8c08b88c",
  1289 => x"08881c0c",
  1290 => x"b88c0855",
  1291 => x"55bf8008",
  1292 => x"802e9838",
  1293 => x"941680e0",
  1294 => x"2d51aaa4",
  1295 => x"2db88c08",
  1296 => x"902b83ff",
  1297 => x"f00a0670",
  1298 => x"16515473",
  1299 => x"881b0c78",
  1300 => x"7a0c7b54",
  1301 => x"a9980481",
  1302 => x"1858bf84",
  1303 => x"087826fe",
  1304 => x"d438bf80",
  1305 => x"08802eae",
  1306 => x"387a51a3",
  1307 => x"f82db88c",
  1308 => x"08b88c08",
  1309 => x"80ffffff",
  1310 => x"f806555b",
  1311 => x"7380ffff",
  1312 => x"fff82e92",
  1313 => x"38b88c08",
  1314 => x"fe05bef8",
  1315 => x"0829bf8c",
  1316 => x"080557a7",
  1317 => x"ab048054",
  1318 => x"73b88c0c",
  1319 => x"02b4050d",
  1320 => x"0402f405",
  1321 => x"0d747008",
  1322 => x"8105710c",
  1323 => x"7008befc",
  1324 => x"08065353",
  1325 => x"718e3888",
  1326 => x"130851a3",
  1327 => x"f82db88c",
  1328 => x"0888140c",
  1329 => x"810bb88c",
  1330 => x"0c028c05",
  1331 => x"0d0402f0",
  1332 => x"050d7588",
  1333 => x"1108fe05",
  1334 => x"bef80829",
  1335 => x"bf8c0811",
  1336 => x"7208befc",
  1337 => x"08060579",
  1338 => x"55535454",
  1339 => x"9bc62d02",
  1340 => x"90050d04",
  1341 => x"02f4050d",
  1342 => x"7470882a",
  1343 => x"83fe8006",
  1344 => x"7072982a",
  1345 => x"0772882b",
  1346 => x"87fc8080",
  1347 => x"0673982b",
  1348 => x"81f00a06",
  1349 => x"71730707",
  1350 => x"b88c0c56",
  1351 => x"51535102",
  1352 => x"8c050d04",
  1353 => x"02f8050d",
  1354 => x"028e0580",
  1355 => x"f52d7488",
  1356 => x"2b077083",
  1357 => x"ffff06b8",
  1358 => x"8c0c5102",
  1359 => x"88050d04",
  1360 => x"02f4050d",
  1361 => x"74767853",
  1362 => x"54528071",
  1363 => x"25973872",
  1364 => x"70810554",
  1365 => x"80f52d72",
  1366 => x"70810554",
  1367 => x"81b72dff",
  1368 => x"115170eb",
  1369 => x"38807281",
  1370 => x"b72d028c",
  1371 => x"050d0402",
  1372 => x"e8050d77",
  1373 => x"56807056",
  1374 => x"54737624",
  1375 => x"b138bf84",
  1376 => x"08742eaa",
  1377 => x"387351a4",
  1378 => x"e62db88c",
  1379 => x"08b88c08",
  1380 => x"09810570",
  1381 => x"b88c0807",
  1382 => x"9f2a7705",
  1383 => x"81175757",
  1384 => x"53537476",
  1385 => x"248838bf",
  1386 => x"84087426",
  1387 => x"d83872b8",
  1388 => x"8c0c0298",
  1389 => x"050d0402",
  1390 => x"f0050db8",
  1391 => x"88081651",
  1392 => x"aaef2db8",
  1393 => x"8c08802e",
  1394 => x"9b388b53",
  1395 => x"b88c0852",
  1396 => x"bcf451aa",
  1397 => x"c02dbfb0",
  1398 => x"08547380",
  1399 => x"2e8638bc",
  1400 => x"f451732d",
  1401 => x"0290050d",
  1402 => x"0402dc05",
  1403 => x"0d80705a",
  1404 => x"5574b888",
  1405 => x"0825af38",
  1406 => x"bf840875",
  1407 => x"2ea83878",
  1408 => x"51a4e62d",
  1409 => x"b88c0809",
  1410 => x"810570b8",
  1411 => x"8c08079f",
  1412 => x"2a760581",
  1413 => x"1b5b5654",
  1414 => x"74b88808",
  1415 => x"258838bf",
  1416 => x"84087926",
  1417 => x"da388055",
  1418 => x"78bf8408",
  1419 => x"2781cd38",
  1420 => x"7851a4e6",
  1421 => x"2db88c08",
  1422 => x"802e81a2",
  1423 => x"38b88c08",
  1424 => x"8b0580f5",
  1425 => x"2d70842a",
  1426 => x"70810677",
  1427 => x"1078842b",
  1428 => x"bcf40b80",
  1429 => x"f52d5c5c",
  1430 => x"53515556",
  1431 => x"73802e80",
  1432 => x"c6387416",
  1433 => x"822bae9f",
  1434 => x"0bb6dc12",
  1435 => x"0c547775",
  1436 => x"3110bfb4",
  1437 => x"11555690",
  1438 => x"74708105",
  1439 => x"5681b72d",
  1440 => x"a07481b7",
  1441 => x"2d7681ff",
  1442 => x"06811658",
  1443 => x"5473802e",
  1444 => x"89389c53",
  1445 => x"bcf452ad",
  1446 => x"a0048b53",
  1447 => x"b88c0852",
  1448 => x"bfb61651",
  1449 => x"add60474",
  1450 => x"16822bab",
  1451 => x"b70bb6dc",
  1452 => x"120c5476",
  1453 => x"81ff0681",
  1454 => x"16585473",
  1455 => x"802e8938",
  1456 => x"9c53bcf4",
  1457 => x"52adce04",
  1458 => x"8b53b88c",
  1459 => x"08527775",
  1460 => x"3110bfb4",
  1461 => x"05517655",
  1462 => x"aac02dad",
  1463 => x"f1047490",
  1464 => x"29753170",
  1465 => x"10bfb405",
  1466 => x"5154b88c",
  1467 => x"087481b7",
  1468 => x"2d811959",
  1469 => x"748b24a2",
  1470 => x"38aca804",
  1471 => x"74902975",
  1472 => x"317010bf",
  1473 => x"b4058c77",
  1474 => x"31575154",
  1475 => x"807481b7",
  1476 => x"2d9e14ff",
  1477 => x"16565474",
  1478 => x"f33802a4",
  1479 => x"050d0402",
  1480 => x"fc050db8",
  1481 => x"88081351",
  1482 => x"aaef2db8",
  1483 => x"8c08802e",
  1484 => x"8838b88c",
  1485 => x"08519da4",
  1486 => x"2d800bb8",
  1487 => x"880cabe9",
  1488 => x"2d8f8b2d",
  1489 => x"0284050d",
  1490 => x"0402fc05",
  1491 => x"0d725170",
  1492 => x"fd2ead38",
  1493 => x"70fd248a",
  1494 => x"3870fc2e",
  1495 => x"80c438af",
  1496 => x"aa0470fe",
  1497 => x"2eb13870",
  1498 => x"ff2e0981",
  1499 => x"06bc38b8",
  1500 => x"88085170",
  1501 => x"802eb338",
  1502 => x"ff11b888",
  1503 => x"0cafaa04",
  1504 => x"b88808f0",
  1505 => x"0570b888",
  1506 => x"0c517080",
  1507 => x"259c3880",
  1508 => x"0bb8880c",
  1509 => x"afaa04b8",
  1510 => x"88088105",
  1511 => x"b8880caf",
  1512 => x"aa04b888",
  1513 => x"089005b8",
  1514 => x"880cabe9",
  1515 => x"2d8f8b2d",
  1516 => x"0284050d",
  1517 => x"0402fc05",
  1518 => x"0d800bb8",
  1519 => x"880cabe9",
  1520 => x"2d8e8f2d",
  1521 => x"b88c08b7",
  1522 => x"f80cb6d4",
  1523 => x"5190a62d",
  1524 => x"0284050d",
  1525 => x"0471bfb0",
  1526 => x"0c040000",
  1527 => x"00ffffff",
  1528 => x"ff00ffff",
  1529 => x"ffff00ff",
  1530 => x"ffffff00",
  1531 => x"4e657074",
  1532 => x"554e4f20",
  1533 => x"534e4553",
  1534 => x"2076302e",
  1535 => x"32000000",
  1536 => x"20202020",
  1537 => x"20202020",
  1538 => x"20202020",
  1539 => x"20202000",
  1540 => x"52657365",
  1541 => x"74000000",
  1542 => x"5363616e",
  1543 => x"6c696e65",
  1544 => x"73000000",
  1545 => x"4a6f7973",
  1546 => x"7469636b",
  1547 => x"20737761",
  1548 => x"70000000",
  1549 => x"50414c00",
  1550 => x"426c656e",
  1551 => x"64000000",
  1552 => x"4c6f6164",
  1553 => x"20524f4d",
  1554 => x"20100000",
  1555 => x"45786974",
  1556 => x"00000000",
  1557 => x"4a6f7920",
  1558 => x"32206275",
  1559 => x"74746f6e",
  1560 => x"206d6170",
  1561 => x"20410000",
  1562 => x"4a6f7920",
  1563 => x"32206275",
  1564 => x"74746f6e",
  1565 => x"206d6170",
  1566 => x"20420000",
  1567 => x"4a6f7920",
  1568 => x"32206275",
  1569 => x"74746f6e",
  1570 => x"206d6170",
  1571 => x"20430000",
  1572 => x"4a6f7920",
  1573 => x"32206275",
  1574 => x"74746f6e",
  1575 => x"206d6170",
  1576 => x"20440000",
  1577 => x"4a6f7920",
  1578 => x"31206275",
  1579 => x"74746f6e",
  1580 => x"206d6170",
  1581 => x"20410000",
  1582 => x"4a6f7920",
  1583 => x"31206275",
  1584 => x"74746f6e",
  1585 => x"206d6170",
  1586 => x"20420000",
  1587 => x"4a6f7920",
  1588 => x"31206275",
  1589 => x"74746f6e",
  1590 => x"206d6170",
  1591 => x"20430000",
  1592 => x"4a6f7920",
  1593 => x"31206275",
  1594 => x"74746f6e",
  1595 => x"206d6170",
  1596 => x"20440000",
  1597 => x"4c6f524f",
  1598 => x"4d206361",
  1599 => x"7274206d",
  1600 => x"61707065",
  1601 => x"72000000",
  1602 => x"4869524f",
  1603 => x"4d206361",
  1604 => x"7274206d",
  1605 => x"61707065",
  1606 => x"72000000",
  1607 => x"45784869",
  1608 => x"526f6d20",
  1609 => x"63617274",
  1610 => x"206d6170",
  1611 => x"70657200",
  1612 => x"524f4d20",
  1613 => x"6c6f6164",
  1614 => x"20666169",
  1615 => x"6c656400",
  1616 => x"4f4b0000",
  1617 => x"496e6974",
  1618 => x"69616c69",
  1619 => x"7a696e67",
  1620 => x"20534420",
  1621 => x"63617264",
  1622 => x"0a000000",
  1623 => x"16200000",
  1624 => x"14200000",
  1625 => x"15200000",
  1626 => x"53442069",
  1627 => x"6e69742e",
  1628 => x"2e2e0a00",
  1629 => x"53442063",
  1630 => x"61726420",
  1631 => x"72657365",
  1632 => x"74206661",
  1633 => x"696c6564",
  1634 => x"210a0000",
  1635 => x"53444843",
  1636 => x"20657272",
  1637 => x"6f72210a",
  1638 => x"00000000",
  1639 => x"57726974",
  1640 => x"65206661",
  1641 => x"696c6564",
  1642 => x"0a000000",
  1643 => x"52656164",
  1644 => x"20666169",
  1645 => x"6c65640a",
  1646 => x"00000000",
  1647 => x"43617264",
  1648 => x"20696e69",
  1649 => x"74206661",
  1650 => x"696c6564",
  1651 => x"0a000000",
  1652 => x"46415431",
  1653 => x"36202020",
  1654 => x"00000000",
  1655 => x"46415433",
  1656 => x"32202020",
  1657 => x"00000000",
  1658 => x"4e6f2070",
  1659 => x"61727469",
  1660 => x"74696f6e",
  1661 => x"20736967",
  1662 => x"0a000000",
  1663 => x"42616420",
  1664 => x"70617274",
  1665 => x"0a000000",
  1666 => x"4261636b",
  1667 => x"00000000",
  1668 => x"00000002",
  1669 => x"00000002",
  1670 => x"000017ec",
  1671 => x"00000000",
  1672 => x"00000002",
  1673 => x"00001800",
  1674 => x"00000000",
  1675 => x"00000002",
  1676 => x"00001810",
  1677 => x"0000034e",
  1678 => x"00000003",
  1679 => x"00001ad0",
  1680 => x"00000003",
  1681 => x"00000001",
  1682 => x"00001818",
  1683 => x"00000000",
  1684 => x"00000001",
  1685 => x"00001824",
  1686 => x"00000001",
  1687 => x"00000003",
  1688 => x"00001ac0",
  1689 => x"00000004",
  1690 => x"00000003",
  1691 => x"00001ab0",
  1692 => x"00000004",
  1693 => x"00000001",
  1694 => x"00001834",
  1695 => x"00000002",
  1696 => x"00000001",
  1697 => x"00001838",
  1698 => x"00000003",
  1699 => x"00000002",
  1700 => x"00001840",
  1701 => x"000017b5",
  1702 => x"00000002",
  1703 => x"0000184c",
  1704 => x"00000729",
  1705 => x"00000000",
  1706 => x"00000000",
  1707 => x"00000000",
  1708 => x"00001854",
  1709 => x"00001868",
  1710 => x"0000187c",
  1711 => x"00001890",
  1712 => x"000018a4",
  1713 => x"000018b8",
  1714 => x"000018cc",
  1715 => x"000018e0",
  1716 => x"000018f4",
  1717 => x"00001908",
  1718 => x"0000191c",
  1719 => x"00000004",
  1720 => x"00001930",
  1721 => x"00001adc",
  1722 => x"00000004",
  1723 => x"00001940",
  1724 => x"00001a14",
  1725 => x"00000000",
  1726 => x"00000000",
  1727 => x"00000000",
  1728 => x"00000000",
  1729 => x"00000000",
  1730 => x"00000000",
  1731 => x"00000000",
  1732 => x"00000000",
  1733 => x"00000000",
  1734 => x"00000000",
  1735 => x"00000000",
  1736 => x"00000000",
  1737 => x"00000000",
  1738 => x"00000000",
  1739 => x"00000000",
  1740 => x"00000000",
  1741 => x"00000000",
  1742 => x"00000000",
  1743 => x"00000000",
  1744 => x"00000000",
  1745 => x"00000000",
  1746 => x"00000000",
  1747 => x"00000000",
  1748 => x"00000000",
  1749 => x"00000002",
  1750 => x"00001fb4",
  1751 => x"000015b7",
  1752 => x"00000002",
  1753 => x"00001fd2",
  1754 => x"000015b7",
  1755 => x"00000002",
  1756 => x"00001ff0",
  1757 => x"000015b7",
  1758 => x"00000002",
  1759 => x"0000200e",
  1760 => x"000015b7",
  1761 => x"00000002",
  1762 => x"0000202c",
  1763 => x"000015b7",
  1764 => x"00000002",
  1765 => x"0000204a",
  1766 => x"000015b7",
  1767 => x"00000002",
  1768 => x"00002068",
  1769 => x"000015b7",
  1770 => x"00000002",
  1771 => x"00002086",
  1772 => x"000015b7",
  1773 => x"00000002",
  1774 => x"000020a4",
  1775 => x"000015b7",
  1776 => x"00000002",
  1777 => x"000020c2",
  1778 => x"000015b7",
  1779 => x"00000002",
  1780 => x"000020e0",
  1781 => x"000015b7",
  1782 => x"00000002",
  1783 => x"000020fe",
  1784 => x"000015b7",
  1785 => x"00000002",
  1786 => x"0000211c",
  1787 => x"000015b7",
  1788 => x"00000004",
  1789 => x"00001a08",
  1790 => x"00000000",
  1791 => x"00000000",
  1792 => x"00000000",
  1793 => x"00001749",
  1794 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

